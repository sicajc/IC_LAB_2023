`ifdef RTL
	`define CYCLE_TIME 2.6
	`define RTL_GATE
`elsif GATE
	`define CYCLE_TIME 2.6
	`define RTL_GATE
`elsif CHIP
    `define CYCLE_TIME 2.6
    `define CHIP_POST 
`elsif POST
    `define CYCLE_TIME 2.6
    `define CHIP_POST 
`endif

`define CYCLE_TIME_DATA 31.7

`ifdef FUNC
`define PAT_NUM 828
`define MAX_WAIT_READY_CYCLE 2000
`endif
`ifdef PERF
`define PAT_NUM 300
`define MAX_WAIT_READY_CYCLE 100000
`endif


`include "../00_TESTBED/MEM_MAP_define.v"
`include "../00_TESTBED/pseudo_DRAM_data.v"
`include "../00_TESTBED/pseudo_DRAM_inst.v"

module PATTERN(
    			clk,
			  rst_n,
		   IO_stall,


         awid_s_inf,
       awaddr_s_inf,
       awsize_s_inf,
      awburst_s_inf,
        awlen_s_inf,
      awvalid_s_inf,
      awready_s_inf,
                    
        wdata_s_inf,
        wlast_s_inf,
       wvalid_s_inf,
       wready_s_inf,
                    
          bid_s_inf,
        bresp_s_inf,
       bvalid_s_inf,
       bready_s_inf,
                    
         arid_s_inf,
       araddr_s_inf,
        arlen_s_inf,
       arsize_s_inf,
      arburst_s_inf,
      arvalid_s_inf,
                    
      arready_s_inf, 
          rid_s_inf,
        rdata_s_inf,
        rresp_s_inf,
        rlast_s_inf,
       rvalid_s_inf,
       rready_s_inf 
    );

//---------------------------------------------------------------------
//   PORT DECLARATION          
//---------------------------------------------------------------------
parameter ID_WIDTH=4, DATA_WIDTH=16, ADDR_WIDTH=32, DRAM_NUMBER=2, WRIT_NUMBER=1;

output reg			  clk,rst_n;
input				IO_stall;

// axi write address channel 
input wire [WRIT_NUMBER * ID_WIDTH-1:0]        awid_s_inf;
input wire [WRIT_NUMBER * ADDR_WIDTH-1:0]    awaddr_s_inf;
input wire [WRIT_NUMBER * 3 -1:0]            awsize_s_inf;
input wire [WRIT_NUMBER * 2 -1:0]           awburst_s_inf;
input wire [WRIT_NUMBER * 7 -1:0]             awlen_s_inf;
input wire [WRIT_NUMBER-1:0]                awvalid_s_inf;
output wire [WRIT_NUMBER-1:0]               awready_s_inf;
// axi write data channel 
input wire [WRIT_NUMBER * DATA_WIDTH-1:0]     wdata_s_inf;
input wire [WRIT_NUMBER-1:0]                  wlast_s_inf;
input wire [WRIT_NUMBER-1:0]                 wvalid_s_inf;
output wire [WRIT_NUMBER-1:0]                wready_s_inf;
// axi write response channel
output wire [WRIT_NUMBER * ID_WIDTH-1:0]         bid_s_inf;
output wire [WRIT_NUMBER * 2 -1:0]             bresp_s_inf;
output wire [WRIT_NUMBER-1:0]             	  bvalid_s_inf;
input wire [WRIT_NUMBER-1:0]                  bready_s_inf;
// -----------------------------
// axi read address channel 
input wire [DRAM_NUMBER * ID_WIDTH-1:0]       arid_s_inf;
input wire [DRAM_NUMBER * ADDR_WIDTH-1:0]   araddr_s_inf;
input wire [DRAM_NUMBER * 7 -1:0]            arlen_s_inf;
input wire [DRAM_NUMBER * 3 -1:0]           arsize_s_inf;
input wire [DRAM_NUMBER * 2 -1:0]          arburst_s_inf;
input wire [DRAM_NUMBER-1:0]               arvalid_s_inf;
output wire [DRAM_NUMBER-1:0]              arready_s_inf;
// -----------------------------
// axi read data channel 
output wire [DRAM_NUMBER * ID_WIDTH-1:0]         rid_s_inf;
output wire [DRAM_NUMBER * DATA_WIDTH-1:0]     rdata_s_inf;
output wire [DRAM_NUMBER * 2 -1:0]             rresp_s_inf;
output wire [DRAM_NUMBER-1:0]                  rlast_s_inf;
output wire [DRAM_NUMBER-1:0]                 rvalid_s_inf;
input wire [DRAM_NUMBER-1:0]                  rready_s_inf;
// -----------------------------

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
as0Rr8SuJLgs/qXZ7YQ2pMO32XASpJEJL7VK1My0LLHVYQZDnwbwGWaJDvQJYsx7
Ekm+2hTPoG31ZFKFBVGcmzqvJCAOuJbOtEU7ojizW7g1Gfm9wbwCITh0Or5D23Jw
AR+HH5p5DpyNzcp7xJuqTkwQjtvuSTM5lPrBwQ6EAds4g3Vkl01vSg==
//pragma protect end_key_block
//pragma protect digest_block
SMS/qnz9qAoTX8SN0GmRhWGwgsY=
//pragma protect end_digest_block
//pragma protect data_block
Ege0gBr4zB7c9I9peye6QdIgPiIK86eUZPz9NeDcLlnKhR0hMqRr4yeuiNB4YGUL
Qzux7inQzF73ranbMjwIQst+lt8td0B/gt3fOZ6qgssHL6+EwWWqGukPtwS8PqSN
9tMo1A1KIyWyEhrPsllqhFscyrBoLTKFxAdGy1DOcoCQYSMlvIuovb4hlMAb2kFS
AAwAfrUa9D39011WivIbOaXofm7CRddrTeiO/z/2D7ybzRCaqKeej4qt3da6nNO1
jEefoDGS69WP4B3e7MWyXgKvN2+IqFLFBHDxl3CAB9tED60iDAfNa//JJWA0HMxV
0JV7ebRpHrtlJRlgVXGZs4eBBHfKfks/7+a8W9uHQ24lF2jB0gnP+ZaJFP39nyVX
Q+AlKIr2XVoDguZNsAK0sGluIsDIstee3LPiDUySi7BYB1WmumwGM3s882ivPEKm
eQjZ1EDUOQyk9UZo+rn8FKCtJJbCrOB6AjmHhZqrQlhhsDAHplEHyw5dJTx3huLF
JkpS3RjZ0iSxmbM5mrsZaqwo6U5J+fveyHJxajVEtkRyuid5A5bhfMME/9nfqTue
gwIBJxbtopAde9jzByhwraWPpmZFch09aoj7z380NfzcrnD5vbZ2M/f0XtgWPcjJ
fNcADmlybDK+mgjDOdDwqTKNnBRhX+AtcmaWq1fybygQIDmAWo0hKNo6OhHhYUe8
Kl4WV1o2ZUEl/EhxO4LeQmGx2ibZJX6OiCGGE60C9u66WEiQmrlBnO4m1aJeG/nf
0qcCYc1Ln5pdhnm3RqONuojpxZgk+hwelgUSfNcTM1m6AjxjNjtwXsA4mQbELL5y
K/nuaw2lsv0NlqSyvCFOQQdWhIArqOglUP0kWDXxaMnbqxJOADwh5UhlRf5PLIux
vDuwSXVPC+EAKqhatKZCxsQGTx//zcL6a0m40fAcwDx/3gUMYCFHwHsXi3w56LAE
4lw0bAA0ua/pvMQLudIwRDB8CBMEKJdxk3MrpPvAOJibhMyo1oisdC22I4cILTwy
zCb15b0ye+Lj3utKIlZaTbEMyhjvdkuDxZKCCQk+BBDICnY8XjtppYQ0vB48IZBy
DNE7XNhwqayen4Ob1zuhnIRKNDCpvsRuBxjXHUuf5kePqGnbbQxpY03kE1iA/y7z
yEn2FlyJAyh9j5eSRgl9mDeUdVLJ8kEgQWQZ/m7RJ2O7kYmaSSansOvHzLKzT4wC
FMQjD0VhZia7Qe2WS5RRI8io6GEaphE1IjjUMLjUVlkMHN/1AWK7ePN3TeFuwYvq
EhRq0lEWsDP/7gVIXVm6kbE3PIdC8xxKy8Bv1XNOxhblpGwPdoixjGe/yywWJXCz
lGzau3rmATmLXx0NUbLcQ6DkU+h3C4kccktFAnlj9MXsa+zSIC5YqF4+Y1FdJGyD
iREwgEoAnePsc0dNbNe5Cx6NQoEazVk+ZeNTzovOAs1QxRLWrtrM/BjIp1iKO4KU
ynbEjZhvNVW8LDwVr2FxIphC80gsfYtlPlNgQ+FdQQE62cKoxSI7Svoc8ukVmk2f
KJpJASes7oo8UmkRZW706iqXmLw44i5go1Po4VudFdDafHiHO2tewXcTqAbqCA/3
+vLQp2iOSJSKLYfWBodii75X4e+31DTxGDtFBa3pNmc09beeKvtw2PX87mNiukti
NZCunJvY+195bLAxJxgKomv2IW+yEB9JJl/+86gahkoJx+hcSN78XCOjRti/dnaR
EyqVtiyDxn5J30bnrijA61FF8DAG9NqglFSJMGnyh8Xi0eN6ZCOh2wk8hjiiE5em
g1ucu6bZTpu44U7uiPtC6vyx0aq1Vl8nwPnoz1uPVv5P4Z+HBcEUPukksCoGnkds
8JDhPjolxcvz56RkF+cDOXTmBklpHaSKFyq/u0GCpSr9R7XNfvlfAdl4kvO1a+os
BaD/57PpQAyLD14ywfjk1jYrZa+pY9fRNzXWsyEAAyfOBly5PrQFg8qbKx5Yu+Ar
GaDwGs08dHlIoyXgrA1C8gyS1caEQUJl7C/e2HwU+nb2s+sQB69YwJhM4a+qpZMY
8W+CeHd3X+HQPPOe4ztDvBjL314RmqVk1xQAs/S4R7ctJ1XUK3MOj14H3rdJSaug
UDZwXWAYVVcHgYt/kaliAgGX06n5aj98EyRzn/JemNXuJG6MFNxKp8ZvICZJUXw7
NLHLGBcf2SUTmRS+LX5HCRm4/VgvpOIgZ8vBP/U+OuOYZ3cs8JiiH/0rAB4L/JWH
4vOmbjMxwjrGhvA9rEeexqO/hu27+a3eQrHL4qdVcoF1EISBjV7V6eKlMwKiyWNF
+eOzB8CrauQqyLHpPkDxLaYVaRxqrk2kyZD7S3xm2/6vL7alrJqymKanLv5fmVCF
gKtGJBMwYtASPFVsXXzrAiZeuHp9ToxEKjbcUYs05V2cnlSmPZNeM/E8xf7RrM1a
prhL2XGNajYrZPencMRohxhXketQBn6Gsnl5eltgciff6a7yhQI33Q/g3MH+fE6m
APRqzVbGymixu3+SB8soVv/oQJlF9IYqF37cuolCsp4nLtEwZRWyRrzWmwr1AcCL
75ORq5X0c1qQkduYLymUMVHXLVJXYnoIa7sF74694eJrovmBicVNNwuXIMO2UpyV
03NREMjPNIQ78nGCZo/A5TO2X5bvMJofxKnEqv7VchU89DeB/6TjWXbkUZ6CJn3Y
LkQfVP5qI7h1lQPL8xXMNE3z1LkEJbJhMEsIljezOAv/EDYzy4r54vauLU2YWlS/
A1RwIw46zDusBNQ9gvgtj/g/HCjb9dNpJuz/LveA/EpqS4a7MIhgc/KnMj0wJD91
YL9tUIa310aqcKkj+nOGbDza+bVfPvc6ImwfaktREgfTcN/4q8m2le6BX41haSoj
52x8fPbhQlD19a9JQVSbOM/lf20NMvQDWZl7H7JzE85y25auLI7wEEOEmLdYyXFG
Ks/fiolIlVNhu34Mlyw3/qSLO9pLbaV9/dxJlfHubwNcpQlFBVuf3mJun+b7PlmB
LSZGKw8fu6+5yvoHCvTbxptHJ6p5XD3u3E2onGiGeuCgzBzPwD2wrkeolnQoJYzf
sdvsMFLJ9O2EQ9+O14jJ343M1OooKfOO8LP8Y5Nh5UFRsIyQ1Hmbnq0oUz1ChQ1f
qdSdqKHpb/q968jFaPNscmNXYtdjbqlJz1bHaHA+e1SiSFSWzW4PSYOT+J4Zeege
PjM36neeOCVGtBZ5VINtY8AYlSm3cH5NPYteVwmhWol57WMwLQWYu4cjVN3RgXk1
60hWB5sA8mmo2bZQJwkAtlbVj6xbl3qEkk3/11aeEiOfF64y5Ng0JpNxX8U8Ko/B
OitKC3F1pcg33pelCse4u5Y0SxE+ZiFmxFqs0MIhvuZhkc3k6z7OMXvIxJE9jnmW
m1/5x63kYiOhHLGJRp3Ji2jRJ3u1AYoEdgATcP6vz/1f68/CpWT7V1koFDXppkpO
LkDddK1wVVQk99hELsrF/dlGe7M2bBzuqPa9r8v7iB0FMpEP3aoQhDtC9AnHPCPV
2xDcWilILe+Zhkzv5cBjiHgRVXsLQQ8RbmwX8bfxJooD2SzpCrLNQjwRRgzMj2Vo
fbXq3HlsGfI3b8Cj7AJQ/AhGnTUGekCC0kZXXd7ArpX1AjDBAvhcqc5ZeCXDdJh8
Tlhr4/K3bqneC4flw846UiTsmiIyw1X1pB38C5FbRDJBQl+vVX8W6dnsW9ON+Axj
fTLEisguqeEu/OnRccv/OADo2r+M1k3TWRQBUHo5nAwSJxCqGMqt1XEdO6ofv6r4
uo21R1vp1rlQD5dZKUHYN4n/POPe3n7Yni79YXB139IeoIE0JKnekjdsTEeSm2Af
7CZHyKODtHBbBEtWTddDaFhvBKcIQT1uoZAkS1/L60I/gPAES6Ke9uIOlhPtlVQC
+y6faQslhzA1XymkbulyD6u+TD2ljRn1Lxwf501/etDJj2bIOEmX1V90IZk2DRXn
zCG2wZnjWM2UR0uf7KHIwsaVqkupFG0gw91gyAJbrznoL8LoiEahvpcRINmlkieO
bn6Y/AVUN4UmeIJd+jMDsfLbNZ/j0iwDFJeq/FqHUesA56Sh2TFxVPa0XzRfNDe5
JG0vD1PniX9Rb7KtQww22eLt9t54kJbibTgjeDvvusOAI7kHVdy9ENpvOVtXB8rr
N66j7IZHMYrJ7yr8T8rHn/0nA53xfLWeAD/SNijLwFFFOqzamq7b5SrDVh14+n+l
ustB/yFvMhdjw+JwA/TRjPQGcaREsGGx3aimy+CNqhA8K/yuzqcAnxM79bu684ZL
5nTgbCmr8BvDiXAwaswSfSX+moTsjPCf5FYo6SsSrsJ71eJCnVyGH34EoxSt2dk0
mGVGYD5Fi6fiSuOYLLqYlr6G8uVOuc6XKlqlYn7Fi/k66yO8jX9PzFeh1GYGFSBT
hGalVAyYUtGHT8gbQvMdntAQyLUKsw6NIpmtRY9JPcqmxj4sK2ozc1mwik9xemhB
AiXkJy7nI+OnS3IYl7GXtduxuN7dYxFk62arHMBHnaPcUVJledqfR5kZF6/e4ef2
/C0SoAIY1fCbs2/Py+K7mjntpqDYk7DnErBtBN2dYgYsfvtyMIYUkE7n2HOawBEk
zDC/IdIj1STt6Fi4m0LfViw6pvtu5dUpkNwsYrlqaKr+0B7PhaglwKalxNNfiidT
MZOgiITSeib0exjpULw9eot31i115DuqbSGwD/P0Ow1MXVtnVcV2rJDPHVP0fTWf
5KFt+Tggp6KRUBHJk1Og+KI60g7FaRv8qgO4Ud//8umAE5wcIh8DMKJlAv9TnIlB
PRN7hmjNgdJIa/1SY4dyPjO2GyGAYnzKVOnJEZFJYqw0m9epUoYP57bgmgR6eLhE
Nj01KpGGBGKXwr15/+oaIi8ZRpKaGZLGrbqQFLm4Ojqd/vDOXVtNS22c3NBIri7I
Uzdm2rXojw54P6eQU7uHsSUVoQ9E1PDbXjEFOpSvcfFt57FTGujidPYK/vvbyaAo
x5KCmPtMArnWneYdEYpEI7pRfYijtMdpMQDa1GcYKRH5OsNqGCmUAzidK+aEacSh
5D111XZ2kCtrJhNb/d6+lq/vokiWUnCjltzRMqvNk2HVMK3ujZSmXPdTpl2gL64Y
pM53qRjN+fVOmFiXxXSB0xBXvBqbY603E6wilc1Oh22VCiZhNCPHUBSiaa3r5DnZ
EMnO4aUHb4jizhI2Q4fMPkewvYFWqPjL0IFxBBySiHpcIlqWihhIapW/W7nQxD5i
FDyxR/GzllrRJFKdfcjX42v5MDvXpvwUy4Ib3ln+yLTvdQ3C2R/DAUq8oVm6M81w
fMbQLJ23TX3OM3gVKS0u5SIX2xCiP/ViI/7pz6uaHAZEA52ay/M2kpvp1YNEfNok
EwJSqxBtPMI1Ee8n7B15vE7ZTWFY5SEdCQAMyARQyc1Ki4g4SyFYt03K+CAHWo02
IlGj4v3CtG9WDiqiIGbnUuTq0mzXZ+7xzHw/Qkf1iE3883+8FytGX0TDLQ/nd3v4
43uO1SUEn79jI/7F634P8DAc5SR4rih+jJN7AGXUPfwTt0oorvxVFSRn32ckHwS1
Bcd1rgIV9EW9oAMEwujQoSm3z4tA33IFpMCoNQAtv6QiXqb8uuDnlabYIXvDJssr
oBdyYTpNnlEF+PIYNGIaceLRxA/eLNVq7UxxHqjeMzWeQSJ34mQFaEh3TVrMnDZE
cb8Y4t1m5Un1EnewP0p6EjTnGFL7sR/a8pFKHSYSs1IenRsgJFdmktQZq4y1rq+w
ZjTULJzTu0SU7wz85r/sYKrDmmW8bOfnD82LszoGD/jYnTNHzZAAo7424Df1POPO
Qery/P98K0azx9CUA01irGKwNE2A3WO8nyFs5FEI5c8fy4bB493WrZheAwvWqnsl
/lQlRupggXaVD844E9Tlx02CwptCRE/07akRcy5m6cBNEfNG/790Gd7E6Jgn2l+p
i3L4W1A+ly83FuzdFe4AWpeyr0a+J4GcQ2AKaBlgckA1cYI7Fh7l3oJb1X5YSxkk
7Tdr3n/f5X26eCfw/kW9YqyMNj0FD15x1soqbXAeBbuBrWLDpoG2UtqhOcE6xiNL
uxehtpt1xQMDx/Dm0qTrdjXPeOEaa1XkU0x7dnP8zUzFqnnPunpexzcbxiOkdKRi
nBM8/47K7hVmMJ5sp3huBhZFtcTnmcgIoxmZo2DbipS8VfeodJatkYYZM0ndBncq
ji4H8IBMgFsZPTyx2/W+owfLZ9kOSNTCaWgWzoeniNFDV0re0fcN7ykd7LoD0wbS
H3RpN9qHj4P1WdqHnMxHPCjmSfKjFzso1tpxi6HIgQWQSHhPdTs9CBm25JSmOTpH
9mmIsm33/tgPeQoNZGoEvOGS7vY4EQHZtoDo22rJeXULMOIjIgvOqQ+tCW1Ed7Nv
DNcy3GTwA7eP/EK0kYrmyVjJ7Tah/l4fxrKqFrcN5CVUjVkDjYd/O+KaL0fn6qra
YB6o8rvPoMwXK9iVGq3U0o2sI0+PAWMKUUCUO8iL7GY12om8yEsMlGjMuEsWTd1e
QyNetKsPXowBGHvMOsHmWHzc58CdkhwZEbm47+jNaExVLUnUR92AjIjTtany22LW
yqLGQFhwqKQ4AG7aqOah+p2QoYKJ85Dp6C1X8qXolszfdICguKsAst0W0a6PT1Ps
ZHCvhOHm0lJ0NvQMq2zED6SuEGErvNiCMXeuzfnKLSyDaAMNn92oPKh5/fM/6tff
KuMqN07HqpMZs6bhROUyGtnCDFcMW9EpinEEq2Fx694pE7Df3/9N8etR7RPobIxb
M1c+weR54EKe9qBNIk1NiP2nMpeSAELeNb+hNx0NsTHmiIUt/Lmn1/j61/G1ynVg
M4FbY/q5VwYcRNYWMK8ma6U/11D5OCYT2TfNkm4p28nr2/z2rs/9XgXVirye+gKE
4xvLankKyM8tYc2blRKgQlzTnE+07U8J6mHNR70rAt94tuUJTWlCO0dTD+eW4QXL
w9EthbOwj9bieLnPaeXnZM7tc/rXYfrn0qGfUGozlZgIDIJv9uFSDHWgN8B5SjNa
q6H/agXCww1u1CQxUDyXRrQUU//sMhhbwdMMiwu6n8Ie02nT3HuAotDQHLuw3iw8
+XwQu5j2ixbX8VQOGjytF1QDP1lF4D2Pmc+tBsAIz9nhP0gZPyRVSlhOqZtqUyAO
8L2GmdQxdwkAiZ+jRy/VoGoqXTeh8WxONmgL9V7UXv9xrhx8MqieOAH4WZ1nOVmf
NRzEYpK3x9/ZKW3eLR7landVBOI/wSku2I9ryRT7aYIZTSD3utwhVvUEUYTaMjD1
1seR9DK6F9TkpAO01Xk+5SuGGBTlsOE5lipXwbN6rW8ERZwELnDAffprmz5fet9t
ZOuw0j0vkzD0HwbXdmVccGAVH7JhGayuHYtYREwTF9k2dk/lV3tFZn2gT7pOJ4nm
huapYqO35JRJG2n5kpYX6KAJVfVkq7y0K+G36dPmXszgPsTQ+M7238Q1H0053VGu
Qy7VWnEhJEY/GHZe2CQFO+lkNNRD/Ts54yElzgfi1YwkHUWINcZBPYifJPky9qyh
kxhjdiSOQqgZKxFkDeXpMet2LZM/t8dJYX2i3VbJfdeauF2tbEU6XhPd/oM77SRv
zNAFC9m8LVFW8gtqhFINsRxQm3Nfrxu3kvH1fWLP+XNJd7MX48xOU7cF/N87hYTA
kz6wIMPNSh80pVhU3vVgfPEodx9/c3EqzRI+Vw2b34TZBjqG/Cw4N1v8/eWlqY2d
kmj4x2F2XvzD1jyUUmnlW6AgbP8us2EGwXJlLYgTC3SBKO7hpuN7TKteQyVrKjnI
IxkWB+7iVl3GU8bQb8i80Xtu5EfxJ/Z1/FKpjD1VrNrF+KBuJFGtG8WdyWHlpLQH
hzvL6zsyCucXVUkA9KLaW2VWqwi01bUpKAafdt44BlueGCZNEtJtAMKfVT0MKDcO
yDVO2dLfBjqHDWRNn8NOT+9tBPzS4lUeFU/JwBaJEiOWwV/BhJT4RPDUvlmYliV/
CN6e3TGYN6OciVIss/3aE7kE5LO1OGjkkjdoXI7zJ1ItCSycfRmHSl8RT86DX1A3
FWEqIZ3uXkOkhMZCMjRachzjGFr8s7LTKaT/VLyWfk3biG/HuenovanPO8A2icR9
+W8wTF+qy7SD0S9CYZMHaIgC54rvz8yEhfgOW0435kgVefrQERLFc+kwbM6EMvCc
F93I0u7wbe54Y+gbUHBUDcRINDUL3adDuDocPZGvAD4edUeeWW7s5Mr1xcr5bW0i
+vtThC/ML0iodV6UkRqXXJD4eEowI/7OfKPkiqZyVR+ZTx+IVATMnk2Tk74wkaep
ZlNFWhTAoEXjCAwxu7C7+13X/+wYNCkgF49R3ju8JdxFVY2UmGD1lbL4wl0Y4Ko8
b5oB3z+1FELyLoIDGQVDbBJJrPP47NiikN/4wSy7ok+MMxrfMzFUT12HS0ac7d80
ETRnEn6FGWCDsiCjZty35EXJwuuff5+p41eHEUgDxbmZEJ58e18rDhRfUkonuiMY
O3vjWZ0tagks73WuDFekDOwvoAl9UecfrETKwl4c/OLTAtsJ3FhwxzG+sLAp7oYB
PHE+j5L8mcME1inHGbZv82QJ67UCiHrvO4g9eomF2PZz5SFn6qFMGpmyNEVnFEg5
nTIMNWAW6eXsAW+QoaC+fPhJrZnJ/9T6h0ICrNUda7w8tfNFCdBXeHX4b8II2H1Q
0H+JmUwbykPrMgXSXr7hHuNZKpdT9jWUyu4FsBbSMk7DEmmFTjkvDM2grIUc96rW
0Km9hWn5ESfD6/bbeF8gp1gooWLcD3M3yFuZcBdyRP8+vI3iW5g/9RndSA3w44WI
+13P+wrxC2DIqtY+Kcf7bd6F7MJFUyWi6w7tPC0OfaCgMc9gV98fJwCHBO0TPWIs
wOS+c/KPDpXnmkui4k5Uhosr8LnVAxS6zWSsIYoZMf/TA7MjB1p/uqWUms6GQZ9t
juHIC/281yFcgmbQJDpVTM79Ra1JT0nlKSMo/SubEk4JNe3EfQnQV2QXUyE7WTtF
0hRYczm76zUwdSRAsrOjSaT8TnnGDzgtAsByFSZ1L7pgFVsfdpVqIlDH0SnDFjyN
NJtQ3LeYUxd/CXSAWH5smAjvMCnO7jhcOvW6k1N7yE3YMxuQBk1kOnms24/GMope
yhuSqNXGI22/ZxvW7WcgNSOEspLnvPCUhll4wXiJYxSjCozsBk8W4yeGgVM2GaUr
q3sn7ek1S02Lg4mOyJURjsS264qM7+W4nGudPiT0iVXn9NcwtlwNFw+ItlNC6pma
LMUlqIl8GBgU88O/kNZ2S5KtttItkYY9xkuiURAO4M8Ah4Kxq7L7HCGjM+qxnv2E
jhbhsemprJomxQ1ZQYrc8JJAdmKR5NcV416MBwM6jr+pb3leZttsq/msOiAShzgn
LgDnDXmgdWEv/0auzY6Bwc02PyGw23Dv7g+VZte1yVFqi6nzBHAWf3YSSmNysP4B
r0XfWOkuh2ZIAgMSbMH54Hn+SU6TKwR++ne+RGELjmOI3Og5lax26IR7jsWdgVKs
dafXRgN+80T0u9mJ+bTtOb1KqMgzUX38zHXTPO4uY8XY+zzWDDJmF8h1OzeFGqgS
eaKqsCcRM1MxddY7h2xm2gtSH7U1tGYef0WhHZGVhCyeuMaAYkNZmjowm4p9XKo5
b9+WgO3dssDkvGKtvaXqgqHCsnGIUxOQ/ZGiUm45tdldUn3qudomDdi+CUfx6XMB
d+2RRRZNxzZPW0gLHqdWOj2BCsO5ruaWaRoZrJRM50Ty5y7def4bH5VgtvxjsBrl
FJqxoCEbOmW8/49YnYhMvwoTDqQmTMh9hzW2D8WGehA+oxILgL/z70N5yN7ajrh2
gQ54bLB/WeGzAGoKTr/8xh1/uE+u8+CK2R5FXxJJRtHFnZ/zuwPoxkgDkx3MWD/Y
K7nbxaWv2gc1ZOXoFJhTPqI5roMn+VhWVynwEfy/XG0zKJiFPkiMAs4IxFum9gSY
ER1BI/0xcG9xCb77r7BamZ6LEevPJ9RmxreksdnbQaexrt22XCSwUVQcLt8fa6Dw
EPqbzKsCHIZkJHtpzEFqgZY1URf5cRlBqdefy6iJpMEmUIC+ByjM60OKtwjR4pAs
2nttZi40Qhh8r3SHJp/hbt4I3npAREgb0E5Piiwv2tWUc68QobRUK0UT5kbcYGo9
XVEoXW0IGtL2gEDdm3U8w7yfQcGygX0XE8f6O3DlvuCFc2Z5Z/XPkVzLzWvk7Twy
Uz8A4k3Q+NWAWq8QsTZz8Keo0MpfgPFELNm1FGPBWFM4XGT0gPDhWx4KqSz6xuEj
X8q13TLvhx6RcUmtzu0VP96pnb9cIh9zL3cEeFEp+knBpSlEfGdoUP7Y3bqDitqL
01HWosHjxf2y1HynrZI5SQiktc0fhzWOancs62gwMhWu3UfF98anQXXcE5WxXqiv
ybgg2RIuaIn7RzawL9pY6ByNtv38udA7g5wJkIWA7pDATaj2NxoyL/7SUvoow9aY
oCY+fgUkxZcUq8JPxr3SNovqT7EiCnGtBgEhtKFZCa4hY6LcGP7QFvtfE32z94/p
fyTfS9pT2ttzK7ABFUGFOXui1lMR9ylmRpa0CyOw7WqenSFzDTqXjaFbxnvXNgg3
bZ2RWX1fRkTRAjbJ7wXY6fOG9Yo1zZjysw8vLxCqn4jabNDerbaOR9kQQYDg63RR
m+vtM72u6AXmXTnWqx34cat+V5dgdjvVwYHDeVdJnTx1q7rq/bIhu4W8cv0wH5k7
21vnYRE9nigKXWC/OuVrY7FWP3CQQF/VGUR9dhNve6LyA55uqUvqAQMKGeXzN7FO
hrFIh7YCWE7D8UgL+igVoaOfP+EzYbnDtsBKOv6GT/CpB8fLtqO05uWAYhe2Uzze
CgPNV8saen2BszQiuCb3PEfOoSjGJLD6Ub4jLSalbvzpRHkcqomVcU8SdHQTVNK5
DTUroG6GkSdmYbBcmu3zFtdilDH5FTBAXGNQhNprNWr3CM0X+QJr9b6R+/5dg7FF
fVfSF0FqbB8HOUvAX8hBqs90yzsFp6Ri6NrDAO/MpGL5j6KlEtLgVIoxI45LWxJv
6yY8WeRR62oOyobp81zcI8CZxO4hJyo5c2cmhpI0fEH1V6YW+UJA6JPtY1oE9WiC
H97r90nz0Qe430FpzSCkX8yy/OOnmMiiNOMxll5DCiLkA4Hs6YhqMme7BawHzF2m
g93jJzPzkIoA0NXXKK+uJxJ2F9w41K2VZaAIsM52K0jCkYHkD9Foys4SciXr1Qbf
GForh8trmeF8duHSonJ55Edz92uUVondxqM8HM7jPhLSIeV9iRS9em0L+kPfzuKK
ZWcLrBh/ssG39o9sW6Nf70qb6+1jjhOQZ9yKBLjKc4mBkF1VeJDvijHARzRPUv3j
mSuXiVQsR0o36ohd/TtjWeIs8vudG1hMf+LTGLfwRJ+l28oehTXQsXStCQeqY3jB
KPhz75f9sCaGtmpN63633SVGSTeqBKqy4GRcPemPKj1SiRbNguD7LuddCTpvWaxS
e6gzkvIyy5maMaKzgIZyyuqOtEObN63VKPTuIiDFpn61CORK6ByfSVPemd/VKbrl
rWg+sEjJ/l47FgT9YiLtwKcJkyUPOTq73RNciidbblSHFlc8Lvy/dB+vDQsVFeVC
0ewFC3T8TXah/3ibcce5usHIIHr8p9mYcdgtcIilp7lvRAJ/H76DMzDunTXY90hj
jzRi05hd1Ji1Uk/52gtYFuuCp0MQKvT8s55D4vxYBch9m4wS6ZbYWo8kL2dgtvgV
g6xUTrrx1QRC/iNzNQogp9gnmYenYJrWUwTphf1rswjSKrY7s3WW7zYXB6tRtnx8
slsDp1Sp/RnzI5967Uhmi48DUIO8KTo50ZT/5JSVtqKPsttrsswO/Rmw463V/gUn
83K40DHRtrCN/MtRk/61U/nngmot4hBUkOhViHbUusVO9RJV4CvSafZZ3isRocrX
k+TVzbRySu5v+99KU4yG9qwtsogwFK0tHV2PWMkXsul4mJV+ZrewDYctOXU2HFot
drrURsuUEwOU178rCmpbZ8oIQM09tbCf1iUN7PU3kbZ6AX2XwtM6T2pHoAbpc5Y6
JCOyp040SLLqacFoJ39wU/QrCIETSscIbFlai7/qUS4dqD9dM+EU5ZcMYQe7UCzh
NRYV2y/AZrC7A1J3HHjIINTa6R0SpQG6C0bQ+uhjSaby8j6P30rElIeuyiAvwGS0
MSIOZ1esIW1n9ZMVKwrJeUN0L2d4Ftl4NvkMreWorPmQYmPP41TAIOY1d2JOfeQC
GlI3ijFY/VmIwmwYA5VAahZrZwBWjpmqXMiG6NZYeJTMrn4Xc7xDGDXBN2jKFKQX
lBZlWTyGSaaRoo3DmlENnt0BDGSRubD3tcpaYN41TzZ9LyV+oZvuRIyp+WaR09TY
Sg21ZcN7kYwgrt4IXowTbXQajMQ0wZg66Y/WLXsAXBn2IKpf5uLFxk/54FdZqosI
IWIPs0sjpCCQfINskrZ/8KhgOySrtLRWsvF8BDkZTM96QUqAAmyHy1IloW+BWRUX
izAi3+RLbNnwCtop8oZQPDjTyJ7YevCpp54YasV/G0vSF6DlWo3He/uXZEbmB9x0
Pcsb5McipuZ2Y+LIn+zgR3NFCrU0N0LapwfnzYxtEyQ0dkx/yaEkbp8922aDjE/c
xu+lVmj618sRVOrMl1dMZtHxWmrQJ9Ex5Jbd0Qe9FAXbPw/Hh8aqYOR0FvKL/F8/
ldhn3QG7iVZIRP7ct0xB/Y9or2UiRAnif7ezg252SDWl4zscAKRoOAt7Rv3Tob0A
S/Gq+eqm5/ZyTsDPpyeFEApgDvunB5t3GOSjzf/N7/Gy+kRIg07QysXxb1onQ8y7
Y9+v+hQcL8QYY6k0nIwuRDPhp8zvokfFecl8l/WShsdcbD2MTiIalvkyuNC6eDew
b4miNBTxru3CjUYPpsEWUI2yDL09Goz7j/73e9ytA8zmBWfSHvTQD725cxhMKYW+
fdwrTnyhc3+yJ6eBHDf08Z6TrUDhw8l//V5Aspx6Gv1Tgo658/KDTTFP0WOHcQrQ
ysS/R94I5eJ9DBpxHaochLD/1VIG9tBCOabvoktzAukJevzWGIGkPaPERG3zCbxS
LB4FTWOTfkiKl9SUbRB51MsPKexfFqPqo2YsAqd6vw6ujhCaj3WW7JXG00KtIAcB
Y/DlfeXjSRMS7WsjyKmnXJsF9WMeFTDIaqx2oI8XIMyFZmfNeALUIfGLuAGHmHXR
cRmPvLKc0x0HppFtsyoOsgwvJTxxdFiz/qjNgvlhWyiOBNz9Kim6f3Tvv06AA98q
q+/uIwwBeid0skGLttK1h8A7FqM2BzZZJFWSBzha3SPXcscxbx5EYWuyB1UE/LOW
R3Lr2/8nabAWXmWUsYetN/aiNWQ7mmVKLxazZrQS2E1mN4rWL+LnrrqiP1N6j9rn
5hWIs5PEkcfcvder7sKACD7lN7g0ZUzuoR9ue6HPu8f6IcIjB8Fp/0qAmKyNHifr
lTmaAXV9xAua0GhawGShCzzsEhq2sRFubeG5TJf3NpM7FKm+l8pmpIjnHoYOwAWc
1myQcpw4rb8Cuh4mSPAK9IxsI0PxrJl6DBvjOJ3rFRXXtKPfxxu2tdpL7MmI5LRf
JxDqWlDJsQW3KCIiCsRXwt9Bvej5HElD7vfUeybZhorE1aU2c+HqJtQ0mY24s7p3
+f/E+JDow+py65AcWwmewU3QdsDBD32d6BU/8embuPtqadvGUHe+t6npMu6JrsIr
YDUT/OHCuGYnCQdqrTg+K2UfqwrWfxn1U+6TB6inZpUiVMug/Sh5EViOPqg7I/13
D47LLLDr3i11/d9YDvxI5A+udnt+Ulxx3NbYmC/LOZLmwHlgD+uR9d6DqmSWrXot
YwnklXj0VqeueCgaqiTrjy/Qo3c7tRyXWx/V45xlYStFHuws4QzPNOXGPLZL842T
F/IDolY+a4dprkZur66Hz6YVJGogZil6QhbRyvgRbR9dr/5AzIymSqW7sNoTz1o3
Pc64czbjWNOcbvSM0qXxSRnC/tdXAsOxD1uvwTu9hMB2I+avCux3JGlebs401YwO
lVLKAv++trUgsW8naaukssac5sDq3TKjUmI86ka2oDwIA5PfpT4J9jkjbpJlrX6l
pyqeRwAkxgByy5vA0ZZrUVCfQ5dYj27mHrEPppaTchTmkj9NaX52/Enp53dXXWq3
mnyzAL2UNDQTQ6wiQl9kZAVsXH1P5dwLG9UJhenaLhl9XNNddgKk/Tj+N0ReMQeM
ktTfPiuDovI5BXG5hdN8ylhZyPCW7AllnNS6cAL6KUWu1UKgv/O689/ikw7hQ76q
QLqHBlHhD6/SYcnuFPP0+BtY8SCNaI9iz6bvM2jYk56x1n1H92wBa9rghHwUl8MP
OQ2juIbYnjmiXphIn5YwdYMAlWPatLs82dDkgir7xZQr41X50Vap/5i1u2C0qqtO
6nS44y6XJyizAiPw1bcIrxjsCkrH+tLaR1+DtB75Y77ri9oXXeAjR7B+wY+evWx6
ywljUbqA3O94Erw4RLKIAl163ce+iQAlFuBT/ZRp64juOtajpZtcKmQLBIBQSUtl
8XukEieRzMra0ScD9vz1eo60BuXQBtSdr/M/Ef+vE2AEjaeKEiKkzQhf+KU3baNP
DliRVolHN62LttMPssfn/gBLKudDi7xPX869xB5oooxM5RkqsXQGDPtU5J0zCsu+
2uZE0bUEkxkbCZ1IoHp4qBqZxvvXKEt2tHxLxPPxpWsxvCD7RfrAXnk3G48EVC1Q
tU4gZlmYZVTB/nP4gEioIluv7yIz/W8LBq7BbH2lCx3+Elll1TBRI2qGgnHPR6+G
kC3F1zOOTpM1H4dscMKAyZdr7RUOeLcjRTlIkW0ZVI2oI/KCm+x27YdCRYqSdbtc
sw+6Ddw1NqlE6e/i06pPVqU4dyUXL1GCWd8pgPLZG6YfQH8tYyWE+n80DhsHsFXn
uoNhLKeYpu80vxzRwdDDXiZCfVD9KbHzm1oT72U6dGT57isDD+ZJYFzYUT4wWNLa
eCyj+LqRzRv44g2y44vle62uKTkPkIW22xOK8xyZTEMsYUHbFEYZMwwiXlY26Aj6
2K5G0N66G1EzsW6j9fOwQ7Y6GlNvux+LWTfG4LjIl2x5SAt5SNAgumR4nUr3qVR9
1otPxXIfcvVeo17hp/4GkGH4t9NOoivtY+X75gjCGnkHG0DjI0UZtkmqAiUe89Jw
HchcvA51mHSpYENFOhzUCV++K57JOPecVHRHYUn/+35kLv1h1Qlr5MtBIAl+hJKe
M6R/5nzNjJRkwtX7C+ZzmKv9Zfu77CcfM8OCFTZP3vxfNxdzDonoVBqcRDflbRoy
DLunn79XHnm10fR5Ovkmwvnb/2k9qxDoAPLzitbHjgxdv4NPasPE8ETqMEudlaJb
MbD7NgQW5avBmPQURY7D8anlnjb2GeDoZD7hiPWC0+FRLDR9n4cZ4hCtFCPy4/J+
trp0OKpcRUGdPskLoav54h09oeRzV3XyNOwGVnoFhhK/gmFpZKlMPRM33/Bj+10I
spEh0hC3Dgae1f8gh5Du0FY7lCJdxIeT/eGJqiG9rp2NIjAI2QNi5eBfQrkskNRa
L3XDnDbmZXA+WdsFbUPn+Et+R7xtUR3n/w2u0cht0aBoczvGIkqqV7/bYKOTKAb1
WohXa4QjbSHvPLxqnQvHZY2q6PkFaVxkJw9VSVwAOalT+EuJv4H/12llyJwwlhxc
oR4EQ75mBrwKX6kj/jbhLlGMfVWJ5dFPdv8nHnwtbQY9mLVflkc39+8NkfX3nF+D
Z36ds3hhN1Tk5zMW1vjDGTFZ+TCqu4wd31oQNFRU+cc0Ajx23gPcXJgDd70TAs99
qpldPK536ZEeSZZJo7NGvGvfWlGqvY2aA8wrwWCIr2LfxrUyG+6X2poXi/vDrk34
NE2cOyn1a5QLUvgTAE8DonrpmlNtSoHm4o5t6FTBgTs17IZUUxrksdWUKpXMM9Hw
kYH5+KwdRGy+jt8rTVYeGeRwHZjNFg2RaHA6NkpzTUe7fvgoNfKbtu5mVx13UNUX
PdKPL9GE6Idl9UTLwWu2WTjtPrdgMGY6BPoUvFYKovtrrOVBIMnHER1bDbo+Gvvj
ogOgwZNh+mdmCnR8OtQTDdGP6BobaS56xGyBX1fN9RP4/j/gelm5ZXCWcBVLwm/n
E1aHo+ys/1vRAnBykv2TbhL/HovhY4NkcPBkTE1QqcdEAxZdjebKcyknoERf6g1+
v8Man+nUkWUUbmYbmGddiXrAZ5qycNj49Hj4rgCq4iVee/1rvCnDx0Bc1jCfkjyJ
VLUFYp5689iXa0MvBtBWnY7lmfKfQ7CZN4VIDZ34coYib1ZfN+vW+OJsJmzRROAl
MZTIoiKvYGlPaI79TzqJtio7i9zxl5TrGAahMb/vm6Zyn5iz/WEhD6ZyR1iOn7SW
MVZVmAzc3BhT+nVTYmuSb3zuWSjiptcPtgHXgeHpFbmDAO2wtuSPn0l+6IrCr/4H
qBuqSCBAYU9DaTt6BS1x+nYNd6TOVzsubP5oqZeXTpTP2HOVcBjd9lZ9O3ADkpZi
IRb+oUlauT0LumRKXjs/6RmTuvgeSFYGFhE59WBTHm9yBRFaxhY447BhkinCJZ0L
rr5HKlKo8jx6ce+LVih20xh9iYl6RxENwS32Nd4Q6pjx1lXLkryO3JO16v0grUmL
eH8pBAfeKsgRTfVp+soEEjdAFyH/5dRRmygfHuR73l0bdNM+VvhJqIboi27Fdjru
bQPr5bsmOfQhVNVqLBBp4vPefZ5uzPbyogcO3J4btRZ0VFEQimaysnEG/MTCLDFz
FPYklI1O4DPU8JjJ1ZCcYEFMwJkAYHgSzoO3oiax58NVdwHFxaSTdBbdw3K6PS6T
PPK8YTcwrcQ6Jr8QZKt9Y74zXKVaWTU5Yn80yRIUaHIFHTZr3HUVzHKVPfUkoJ29
GDzzOOIRPZ0lnmYV+tkIHsbvKEygrEYqdHPppDuiz1lbQscMJfF01ecaJV8gIRkN
3AKnwHhppsC1oJR/VUqv+KJo+PEpm2mTJ5SGh9gZIyNMx31+m8RExumi9vbgc+Nz
pmgwIGN7Ue7eQImk8V9BpmhTLI2PGE7qENnm9eK/qicDTtE6lU97cCZtISyoZ79t
9hIMOuFahgNJ3kRy6Ua14Fw/HrWnwUXPl8bWoGP1OejCPdYV/iRjx3F07BpPTbUT
B8rmvqKUz+nNMRulrBV179BQYgWyp+gGUe4zZ7K0HqMRpsBDxiGMgpzppyLf9yll
W6UbsAPbJRwHTE0dNxtdU2ltaLhJdrQxUqWW6d5LK0XkubPGMDBFZi/OTb3AIKT+
R5UPJjuD3DV8gWsI+JI0rXUz9Rp9uc45qUNF/F2n5PDhu+pa74MBvpr2Mk4FPL3O
F1JJocVkTJl6zAVpnjc1iY0yaw6vnSgAr7cPySRZ076VHtBTUH7hKhLBvYOWPdpK
4le9n8B+9Lv4bRfrNSjzn6NTt0gBxv0r2BQwxEXc0F+bnUI+HewsqNe8rS9JT5sv
1C1H4ctUFNyQ80bi6nDqeqtG4dOW2xsfq//7TRhXX/35AMilctTGX78V1BGAlyvv
OHvFOYAjVAKBTW6hDkJ3KV7s9sICoyuXlJ1v49z46ll8U6NVNm4pbRJ0BY7S0bgI
SxVazERiv/MYO4K+0O1uzkH2WHGwWrPcEfFg7W02+p22gpeNmUspHpt7KPD0tOFR
vL11YuG0f8qaS4J4lDA9C5j3EQLm0fZzqoBxN13tX+mMRKt4RtZuhRhBFrrm/OtO
cpAi89ch1/5F3EFyDeqeSMwxNi56IBHHlvIpkgmMVeaBib4lVGxpVGf1VR4/2DiE
8m1x4y51o0z5Ro0SJfyXc+SRqpsuMjUR/BogEKsTOGyAFBZD7DvYYkj38To/OZwF
0PSwXtb0bRlwI4Hnn/zIfSt8YlK+4Bq9d/lTFxUBKoFriM41S/LD94fW984bNYdW
AXZFQpnrCDT2tGSYDXuWgTNcp2/DNPV0kOTqqC27gqa/UeVY1c3P1fm/o7sw/3bz
OUBTBhr2N+iiynaiZy2V0vVW/Gpnb7VqNOxUUXeF2JGf6lr0+mjNMjqpzhZni2QW
sIxPPv5Fo5T++m/2JP2sQipJiFPW/wADBJNdNmlVe3A0jNd6NbugKkROSVxv3dlv
guQTIXbfco28bmlQvLKGL5Jwzl7SfNKcP5YzZtZcYDqUPmk2OqwT/dYpx6l/HsNn
gy0Fh+y6Rmy/Wyynh3xdtqiAtqZEnV97CseflwBYEb94UkddLKR4k/d6nHSd8lQs
rHLVRhxCNMOSc9mAYxddNA5mojDcxJJUul1JBMfIp+uC93O3lnakLitC1aznsRHl
pP2GC0JVOQifNNRPwOuAIh07/o81pe7M8UskY8tWR7USgoJmuTA0l5nmpgb204bA
57lJzSrwDTxP2j4txRcQjBsn6/HY3kjk2xKx7xWe4UA8Yie0FS4LxK8bfZRWA497
Fyl0oNLFCXpCdFLUR5ea8WfNh4BNSCg28CiIoM5RDU1DICjnXSjOBUfOlHISMfPu
xp3qLoia/Y2m6cpGuKD6vjwz23A0qC3THEffBPZZMOegIA9UFWC3n8u9KSFM79TV
O/1o7QHHWaOYZXFuuSfgPjcHYFnUJkFjlm9nSeEk2zvR5ngu9n743cPXi2Dz6JKM
WFesVTo7bVv+LPB1Z4s0QdzxxHtOt1RbguNCZ1/jv8S8NjXLCMeBKFHXZ6VufwtR
19AAL446RiMDRuSttWR4jnXVqB27EEZKwLDrkXSJvQqwIgML3s3LQBYmkIC/xaEr
gdoc6Mia0WabQ23YMaTZdA9u7A4KuxdrHmKNd8wXsaQU1D/j/YtSEzA2TftGbDIu
oTSSHwRQ6H+EOts/sX//pRHyPyFMKfW85BHoAeJ9rlolCSZt0gmICa4rayvVvO5W
b/IBQuXrJPd7NJoaZBuHDskkrTGDqWg9gMRaDV2jBvdBk71VQyZLr4tSn+Z6d/lQ
zEVl642BDxuHLN1DrT1u6I5dzD5s9oXEHwUQZD7B1IrRKbd2wfc4HoBzpgnSOQgs
pXDUvZ8+96c1b4S2Dw5U+7MP3Y2iQZv2RA2+sopZFntP02SzNGDI23lYNdu+Y8AX
fvIKhsMFvS08xYrSroBlniB1FPXhx2Qpmz3XTu4lL2u+ocN3f0hLdlIs3a4qhHF2
/cXmrsc0UaFExnO6oQo7ZyoL90AWzXacSxicVuZzoDkMJnUITJpCzDqNJwoJ8L+L
hj3K1iG5wP85JrnacuxnPxt77Cr80km98nkLlXJiks1+bopZgM5WuUq7sCQrhZf+
/HBmMHfyc4lGq/PzBzGDuk1s+GuJvSxTyDYz53o9ekUAf5ERu9P6M29PvIciHM3j
6Bf3vY29Lm31geqJCpdOL58lME0UcaU9Uiu7fsf3mIOIqioftoQlnlRGb+ItqG4X
Q5hAziQKprL+9trh7c03P184vvosmGgpmUeVrboolCKn3fFI4E2Xuvyu6QcpSWV4
zaoRe8Ea3Dgslgq+hDNY/T80+H+mP2dTYZYWD/Rv8wRIbmKshOgqMJc7BH41yq/7
aahMTvqPNLe0oxRxUFlKzibgYFVv9fNRLU9qcXLxIUg=
//pragma protect end_data_block
//pragma protect digest_block
LU0AnbKZjJl3Nk3r6G5ssEQDIYg=
//pragma protect end_digest_block
//pragma protect end_protected
