`ifdef RTL
    `define CYCLE_TIME 40.0
`endif
`ifdef GATE
    `define CYCLE_TIME 40.0
`endif

// `define RTL

`include "../00_TESTBED/pseudo_DRAM.v"
`include "../00_TESTBED/pseudo_SD.v"

module PATTERN(
           // Input Signals
           clk,
           rst_n,
           in_valid,
           direction,
           addr_dram,
           addr_sd,
           // Output Signals
           out_valid,
           out_data,
           // DRAM Signals
           AR_VALID, AR_ADDR, R_READY, AW_VALID, AW_ADDR, W_VALID, W_DATA, B_READY,
           AR_READY, R_VALID, R_RESP, R_DATA, AW_READY, W_READY, B_VALID, B_RESP,
           // SD Signals
           MISO,
           MOSI
       );


`protected
IF\3KOLA\J[HQ4-+4ae^KD6e>)0GZ)TN2DH_AETMGZL6b/+I#82c0)()1J#ff?<3
DRO9MY3,?&WROF]]GU)TcDaO<YVD1ZXB@$
`endprotected
output reg        clk, rst_n;
output reg        in_valid;
output reg        direction;
output reg [12:0] addr_dram;
output reg [15:0] addr_sd;


`protected
SYWFK0,2.M4EE951S]gF)QF0T.DdH)bcO)D[9f[072bIK4,F#A0)-)LU@(AUOE&1
:U\Z2JJV2d9PeD+4OO_[5RS-^ROT)-M\L5/-<QUKKGgIB$
`endprotected
input        out_valid;
input  [7:0] out_data;


`protected
;#LfDg#VBUFb=6.TW=7[;YSU(I-&G&bLKWceDC?g+LM\BW5C^+BP)),BZ5APC)1;
Z@4g.^I\:=]dBJGGS4aP8_>):N&5aUF+UR5Z?d-+g^38V-9N7KXS^UIKT#K\1B<<S$
`endprotected
input [31:0] AW_ADDR;
input AW_VALID;
output AW_READY;

`protected
J8WgR-WCd&Z4U8\K87AGe<Ha(I0WN\PZS5\2W]\;,0Ka.#/I0WVZ7)[^NE+6Qd>V
;7;W?QB\NU7]>URf2BaR85d5141QG>+3?$
`endprotected
input W_VALID;
input [63:0] W_DATA;
output W_READY;

`protected
)Ca0Y73CPS89BGT-2Z[OKV:_O>&CM?d6R5A8.D=NJ1O_7GT9VR8D-)GR@W9FP=fX
2T3]3T8OeO[;CZ>F>,J#<C@J]E8[BSO.ffFf:@@URd-_C$
`endprotected
output B_VALID;
output [1:0] B_RESP;
input B_READY;

`protected
e+(f,a928#e/[-;B9TDL90A878Y9d5CY5#1)E>Fg4.KLd[0904eU-)5/c+#JSO(b
DcD>82A#F_8M)YJ?fZ=GLDZ53K/-P(g))Z7bZSGb4FFLA$
`endprotected
input [31:0] AR_ADDR;
input AR_VALID;
output AR_READY;

`protected
HCg<W.R,0e997#QV-^VAN0MS<-/Z9#Xg.g[^&IC^7D89[:S2D\<6&)0E#4d4-M-X
#?5S1KEM5V-CMI:^49H5AA/OaG1IN+gP>$
`endprotected
output [63:0] R_DATA;
output R_VALID;
output [1:0] R_RESP;
input R_READY;


`protected
A)0eFZe8M4QB-^I\dTc-KY+Cf99S0.VZ/KcV2WGZ,F8g3Fd5+Z7Y))LC107?34g@
,6>)T?)6Y=3;b-S874:,[)+C7$
`endprotected
output MISO;
input MOSI;


`protected
QR[cfR;4I.X:UXNY;K-FOFA5ZA<c9=PFKWXUP-cT>F;9[Q3_PQLE3)NZQG1^ceN6
gM<^#3\ceJB2;=45#^#_18ZNT6.<Y(1;<^C)EC.T[>DM0##^Q?VB=W9\D=aX4F0<
5@\SHEc6X&ca=X(3-_E,QES].,KZ+&HR9.aJb,[b:U]M#,d#dZH3WS<Y8bbD?d0C
<7#aHZ(F/AP/T>T\YU?M(X.=YAd:M9N:9Q;-3^^T#R9)8WVC2D>YWKJ7CZZZ&cA1
S5G/5C7PETMW\Bf-2>3@[X@-2EV\D\YIa,WcMY@B)ZI]Q_a2WOF^:[&ZN2bdX;_.
,(9X\S@_^I&f3.7U)d9(fCHbX(A>S(/fV]D.:C08O#9[a,[7UZU(:TGFX^4_ZK#W
5cRUceR_IUE^7E/W?5H5N0;ZU:M&cgNKU0HEFN4Kec.,;g/W^WWb[F2>\6&E;AB8
DFD_1X?I?UW&/E?H3HWN(aV^=[P9&#(dNWg\^_f#,S5.B9=7&FIN5@TVORcG91=O
IX0TdTJFR-:/_1a7BQA=2BO9QfTIT#MKcD<Idd9UHg.0;XF/9:IRdH8(e<^>;W]0
Bg=Bg]7Dg,O.+5469_bgWbe-#6DUE5=)8KVL]Y]_YYKUM##,KW)J[E9Og.Mg(eAN
:H(GWSLMR/AGH?U=6bD_3H7b,XMIMUUS,4F7UAW_H3,\96gMLWXGbT5d-(S#INKT
3-7QHKAXR2;=>LY;.A:1=E<4QKbb:>N;Afbg6>@7gZM#,^RBa_EBD^-EF2;@>9PE
>/LSeW3P<5W,&8eM/.Z[bCRS1fI^cD_a<_8d?+W;<Gd7Je^F6?GF;UF(]AXP1V5K
Ee^O4G\D\E2<:UW3J8U)@)2ELA=7:Zg69<DfU7T)f58ACUcLgKdf9).#J\/@,RBW
5)cJN)Z]N-1.M3-a#/>BC;MJT&1Q>;N1N=[Z88AP^b0./R[=La,X:HbWGf#ag>LP
@/NB/#O&S>=WLZ+U604/Q,_2.M8H<\QP5(GE=T-IDXNQV:7UT&8Wd<F\.HTO9B,W
[#M+c=PNM4aV#dK&5:eeJ\>[J4?;Y9CLgVW5NY&]g-(S8aU\/411gca(02CN((X-
3L#=SZG<+]@7(-X]7QdEXDG<_A=RA0<f]Pa]3&K,5SYU+)1HAW=7eVJK9ZJ&[21:
;5dTEN4d7;\FU2+P:Hg/MRf1NE,N5S41QI,L<(6BM<HCNEeW7MHQS<T2-H0(+Y)V
?LK>-#UF[WZ&RF>-W7YOS4@)MA91=(B3GV0+0,AEOWEA#\XA7KUGEg^K/A@;@WEc
YK(NYf+]AG<f?Q.)U+^#C-76<[D+d3I:&79.OE3ILSa?I(f-#2_E1C4DLUO_NNFU
]]#W?8RR0)073d;68^R=YH/0BEC/]FC3<[=WbBSBGTC(.g>R.L1b].a@^c2>&dVf
;KWR3Bd9OB8:A4YSIgE;@G[XB@^>YS/DT1WR@@8?g/>6PAMI;^?b>=-S#e24TGf1
LBeP/O-\_-D?&77KBfBWS@.0#G&^,@;=60&=aaVY,2N16@ae;TI=F-3YM<FdB=?:
SENMg-7S^3Xa9];c:#CMF\=Z;(?)=Q910M61N^XHf4&_:H786TH(P6)cLE)CJL:1
cGSaM+#:1ec5IE.V9^JD47Wg6WI?>E081W(@\/X0NNbQa<Rb-H,-2NIS^Vf-T<[P
5Wg+29E7PGT_1=<\DJ?LQ3K,8&5/5fdS5RaebcO=1@1PY5ZFb;NI;Ac2b7#UO\RE
P;P<1A->YcM(\=G],M(0g^MZaTT(G[dCJMRK;g>c#09M,WBMA5@GZS]9,S]E-[]R
8ecS>gcFX4?YX8[S33fMM9((+>a]Z+]>c0B.Ed[0W=Ob@W-Y<V7/Z2Dg6(-3/[;9
]<2&I\?Z=c6WKI6/9>>RA[XV1GK\1FPE/3daCZ##V?^&@>)I--1ae?L?-#<ZSW:A
[GZ@,WP<[E1N<>EA0\ZE3EGJOHI;d76_fBM\E-S0(M0J]_QC\#NSTW\86a]X.(fQ
Vbb(.Z(,G1&N_,\6;]I<>=5#IJ;/DN/ZGYO&H^7K?=J5cM69#bG>&DM:?gf3S7#R
9J?Q?BgFg)(5=Hg7eV,AOG#-WbI;Gdg@]Sg/;cJE];[&YbUA=?RebA^FJ)5EZDJ(
88\d>a6U[EY3bA:L[@:cEY@@8M^aBG.E<2NLW?N.I)<\J\QZ9f#5A@W]T55WJ0\+
Ud6..SE:>-V/#Cc8C82M_D&6(;QX=G(;\3,FYAA;Vf:^7AQ8I=:4F3^:d1aV&Y3b
2#21_0P,_(7KdH=bVbG#c;=:99E774OLg-6[fO(1?LGfL?QDF17f6)DK-.V_D\&V
ZN=([\)..T260=GQ5GV3FH/9H8)ccJJ.??OJIA528N96&TW7=N_OTfa30aSL7S-B
FX[F2UQ9GO-/[f,7bCQ7AVV8UX[f_+#&-BUL=4A:<^^8C_+EaBaY[f<Q3b8N^;2+
EHL_:62D8<FEZP>LN.X9MY<XI0[=B>>_SaF.+-5I2I>)LNCb5]D6O-.28PbdMZXV
9#fJ/6ED)C.4-]Eg]d0bZ(+<OXNa89J?7;LOO._7QY:L+04G=5L5cDZM3Pc,OLXd
UOFgT3EEA[Yd[A7Z=5>5N4+VRQJ=SPCTD(a93/D=_E:3_Jd4AT9KL(b,cEB^&4DS
DND;XE6S2=,54FUaSAD3SAJ<6EKH,>2Zff17+&IM[,N+@SR_9_.]+02EgB0QdR5N
Kd8G7&R9B_NGOc^9g13;Y=\HKT2=6F6HAG\dH8Ca4AJO6;G_5ASFF-W9BZ#+Zf(\
WX@4c.((;]AR>KEJ]>+@2ZG57FgUcYH52294>JP39d\D0e<bbQ#UWRRdD5EQC)eI
HT5Q2FYR9CAW]A5K>U\5DdV].RZH3-;/^#D(WPG899g-AP81KSCV-R-RIL7AM(&Q
Nf5N,H9I05d5D#fd=Y/Ub+U1@R#WU9S3QIE50]USf?c5:MXS.E=[JFQQcV4S3;BJ
e-Y)^K#^M4bce0-e?2G+392LJ>dSCWS3a,(R[.bXFUZ.]74.8CB(3U);?_9f1;Y<
1^e?dORKT>\cO?/c+3A_O7XPXE)T3F3=-_F:,#D508M@LVZ.8d3P>gE_#-gc/OAd
L_fUT#DCW?[6;LbedRLNPPeI(1:VLXBOQ#+K/1Wg_@#&P]4D_,a=\H=G</T:gS_5
,MHMeP81d:2YD:f4]VF^]F:C#6.B,TSQc99+L7Q\[YIES[(^HRQ9.(fPT7\;4[:H
G80LE\S8SHV8(gI/bXLc<A0?1>5H0Ce:VN:)XJ8NK)Q5A0ABQN<]X(ec;X]c+fSV
O09O)SU.L4A\S//8;.K[&=:WF=XE:7_UYEC4bAVQa.S66_6W@K5Ldcb_@10?<6KU
.M?=4Fg)>VTc:)a#;4J]#^U;JHK;H<B\>c,@6+0+RcR/4H\G34<GDURRN];SgOXC
;DEQ?IC&G[_MC.=[Z^7#46FZ9P/L-J51B.bR+7O+9A2JNL):OZ.3HE0Td.,H,8>\
FU:KI6W>BEL=S37LNfZ7gQBaG0#^ULWVS1MgcWP;>W/C#0_Ob38))/#c;Y52-8cA
0A/>EOA:OS6KNL,3HZ)=)RUAV(SYYAKb\N#_L+FHF_.>NFE^MWS:CT1G\ZZ3d/0R
6_-(SHRFTQ>BaV_QL/S(-^cd1HD.b[R\&<DQTH.H73#ONdKRBCdd71PSXLBGK2RW
aD3]&ZfbEWd<E2B[G19WScYWe_^:?cAAMWD(&XWB=W[ZT@YGF6Nc&)C2(([RISfC
/H17QO099@THYT3I2:/)PgYc#eK3_b@Q<F((Eeg.1)V9F\ed8=RL:QTRX<U-]H3R
805ZQPc7-e5WT<26TK<G917<0K=eZ8^HB3;-HQ2++\HgG=VI4<-EL;Aa(HO--&OI
O+B-)T[)..F:Z3a)KV:=[XW)ALJ-IR.cD;E7SdY,27?@ca.:0Ya]#)T64\3(e<_Z
0@<gSYg&_Gf3Mbb)Z76d@7Y.KW0]JW^LE>3Y<1T4SZOcbN&?g)XIc+K@X^^@JeeP
RE,M,JEMW8B4#LA>f);5_bF6A<1]:RA[aPMD&E6N9bD/WF,.)2>Ce+CIVG0]WNb2
fBEVVF.b9f4VHZR5;].Y(>;.ES0Mce7-:)9QE:2NZAK3KP]M8E^X>Z;(A/7>.XDc
[>d]D[-&6,5YZ.^Ea>8TME:9]FY[OM5/P2(\)DI#_L5[0@Z\?;_fKKSd^V95\IZS
<@>9O,/SWW]7LI@ZeW=T5PaH?UI(1/,K8MXgBI99I;]+0CA2,]LEH,RK0F#JR2:T
&&9?@O)Z0e:^O?];Qb<OK4PEC^T_ZQ4B9_bRD+R60ZW#G/(ZP_65Q&X@WTO;&,1d
aIN8350I.E@N&73.&_^QU4P+5+0O-&I?#N+L93cgf)=?)+eVW,>^Q&859C[/0?0R
FHI0Ma]d8/UP)E8JE6Y.Cc/59>EPL.cfO3dN.N:YIISSG^?L\gQMZ#LPcfbL8C)@
PL[V-Z_UNA6^bOKCRQ\=I7SP[RAMIABDfO[LLWE9RG>gN?@S5c76R4U_RPg2Y>f7
)SYYMgFCb+0#WfT@Of-/=7\bfNU;TNc2#fV(E@Vg34Jg2TO8N<2)M[4CAP8+#cU-
V:T]B+a,9JDKG&CITPKI3E/(MG#QHR;\CW=PXC54)DX+D)#_&J7#0]BW;L8/>Nc0
e<G@AMGE\Q.,7E28C&dEaKeZ3IdHCZ=dXLPdNIY04V((BeD5^C\6d<(^Ub-.27[P
]5RI1A7<)8?/O//J@,aG?SYc@Sa@U7R\>R1(<f1NdPBbT\NR99L/,&&24cV9=55,
Cg7:>Fd?ddH04.6IC23-NUV].;;d0W]fYSN&,Q6Xa,8)NU?53@0,fQ<[9Le(LF)\
FO,V8()5RK8,W7[&E)4]<4<&WMWQ#Wca1?,48U<d<\QS.>JNK;f(fecefC7=57@?
,Wgd>d-VT=OD+g57O<:Z1+/Z/b7@OH;)ePZ?ZPS/AZJ>SVC8)&6-4MKBB?ReaKKB
&6,?,NV-Z9;NWNJJ=7#84<IJ./5-d]g_<M.H:7;PLA6fUF]VMBA=#XZd]g,Z7G]@
[22-73.O4TZ,0f;9d:\4]7T(f]C)OG<eLLJ=;+YN]8@?(bZgd-D>b>:QDZg\(UT?
R-CQ6DG.(SK\N7@c;F-D#DLXY=#1,EAU<1#@d-#.QNO+O[-C?bJJ7#5G<GCM<=&S
\0&Aa-2F0@TS;MZ<_?Gd+6FVE]7T_,f.6LR0g0&8>NEeW[AJ1-B^R8:[L)]6HEd/
^73#D#7Ga0I;\&A]&dS77aQVZ@JOdJ2JG32Q3\\6a=QUd^:d;<Y&@A@)]EXf_=66
C&J?:FNZDT925f/Y>O_CD9f+X^BX)Ze-]^fBc=cDAT8WO>CHUOYA9T\<EYUN1,?#
gH-#VfW[_CCHgS_M8L(/.7LPBR[TT42M@49<D.bT.6R;ca7T^KXE@MR6^3Sf4KB^
98_28eD0B>KRcL&&Yg=FA?Z-@MH6H=b;F>T>7:#\R2?>AG><a0>A/46M3T.][_<W
XfP+Y3\](KS=@a7UQ7F;^VSRU\ca^TWgC;G4TZWa.Z]<Ga4fRLS@CZ+)JVTI8VR=
(8;Xc)g,QIMKQQ#BaM1.Zaf0\N]])c[ES&#.H>)#Tb^1#gO38gOaJ1B&ZgWV;fF:
f.(@:O[g^bb:aR&0YE_b@#/d.)f(@[1-CfV_3dRMZDMZb_cQB@Z&)G_aAAM/&+)+
@U_gUW_A.WX2[WR?>/^/.0OddZ=Ea1<<A-UgCF=/(^aG,PJGJggGJ558D_YT(5Fb
K._YY3cCM(SJP?HGM2,36-^)_NAfEU:4(&BVUTS/RX\^JFMTU02X:F+&BB.8J=G6
.CKc=8YVdLK#GD^>>@F_C^fR?QG==Aa)L&=FS7Y4B3+)X&O0ReF;_cV&d_WE>E[=
a<2IJ\Hc(a(TS>@<I_LPDZUJ<LJANP)Kc#>D_6?;8B@?H@D,8=Y0g)b]cI99gQ>8
7Ybc=)#5/U@R3M0_[LJ3KUa50WG^DE9cI,bN/:/#=N6LG&SG>UBaU3\TOCa-P)U@
?Y[O7S?PJ_TU::L=G1E32cZJYc-.a5.=(Z1Gb4f>fN\IL#-)>,U3ZcGEO4@Y]f#?
018V:KU\bDbg>T&R/&E1FNa9g4+5\G>V/EYQc^5ZW#(,RVIf3ZZf?;0DS.G6=<VQ
0a-Y;^6:S@CLDa^H^0b(SV@(FXdIe\WB,B,9C1+3,OfM8f\LW9L@UI[ag5>[EgVW
f:Zf5\Q8^Aa::FB)gR>RfE/d+B#9/3SY]Zd(C5/Xa.gA-8ZU92E)W]QR>OCSHeRB
7\8Q0P_Y>-Z<.=/]Z_/<3W/G9J>[OafW.NR5C=ETa&OS0#>-.KPc&e88B0V]FF>H
LbY;F6c1IDICD@P@#K;WON?GV.C89+H/5(9bO1_;@FM943IP^A&aNK+W0dM7@^;+
@(Z^BFX]]Y#W3(Z1X4g8J<bReU;3Ad=N/B1J@5WGMF-?^1)XF/NUa&2\).SF6_E?
GF:#R#20[VT&PQf.\Qb?/R1AN;[a\eagP9T\fQ?^:c?_MedcUCP6gD:STNCb;W?f
0+>EZe5K.CR-)@4WU&(HGAXA3ZM]2SZ\YE_a[]@V.D)f0NHY>dN8;aRTT]fC(0UK
9/=YN.<=4e^AcS;K8GA[10]Q_>AFF<Hb&_a\.HbbFLVA]X#>d]&TF>;H,eHf-725
PO&YN)4VWbM@?>^89cS]Sb7f#IXO;)\M(gSKQ5-O5?@2MXK?gdN,6M_5:7RZ^9Ve
Q?HV,B=g12T@XaMBS19(XY_VcZ6\L<dF#@CZP?Bf2Q0CQ5\Qbc-DJfK:J0#VV[:6
=;<N+E=Y8+22\DJgK-^UJPV@E\6g7X<-(MUKU@,R87E-B;bHIgRDQ7ZcT,FNAPGa
aVAS8g&?:^E<Ze8J]](\]59JeW?Y07J9_I@Bc/<c5[TLGFQJM2>OEMdMgQ-ROC,J
gaTFFPXL_fR:TVfc)KNMJGQ3TK9?:;6P/DfHIB)W=A0KL+SJY&.<:;2DgTWZ.>>Y
>[OD9OHH:-P7^OGZT\-Ob@_+V21W@]_bPZ)#7[7UHe?874Fa@X\OLQIf,VU3.Q_.
.V_03:>H>I5GdJ1XT/FW.7e\ML>K_0H#EMe)<=@;CF7aIOS4.34,)>Gf\S+;R,1)
dX.LDS[L?)=6/gfNGIg#TX@XQ2g>BW\8.\CU?/E8?.&&I52A(JW--P[:BS5Y,@Q:
cYP7<6MA83agMUcAL/\?W=Yg#]3R9Z?bB5B;P98Ec<;97[3QeaC[+V,6X[AG?NTR
&^+3)Tb7CS+ad9#c/II)2?RTA;RCgfb6U0Y4ZX2T[H]+]Mec@DMU1A.C+JL&;df,
,;,=CCJTfVCA+RC9UN&VMX8TP53L[ZH\/_K>1I,CENH^S]c7G^+WMd-3R1K0,ME1
3Mb:O&IP+UcEgB\Cd4^BU)e3&bX)-)e^&9<7,3&DN_Ve&b=,Fba/N++Z<71fVAU(
G+a=PBM:Uc?^W.3;gH62ERADI,E=GFCefdYaeMcffQE=Fe]=_T/VfbA@287[W6(>
>3A\0ccT&?LJg7AL:F]PR_L./4UEWcP0#Z-O;.P?VAZcb[#f15-?&OGD[[Ug#KV;
OQK@RTKL7JA2;fLJ0LCcA_Vb+,O;;MIcXgJB1I(9U\0O(C.e/A;Z27@a0J<TI803
;^:S@1ZA-H1RKH/J7FAcLS#>0_R._YQb]MJ(@BR)?1ALBZWDG<1>S8>S>3P8E&XE
JOFbD@UW=f>/)^gK>N._7M&<B2YJM5K92CGNOXf:S/Y<RR[?DMc.+W(9?QSW/FMf
HVRc)_<=CGbbV;;R\JFNgYQ)<22-4HF4#VFF8IO[/91a&D^^P@@4A1&dL&&1Q_IQ
;F,G3;MI@_#d#N4:8ZbcMb(2)]aJ]0g4=e-OA(2eM#W5YUITF<A4DPgH6gV^1U?6
W^LBKE+\YU4\^/N,&&0LQO,-1>:bLHb4=9S:F>-UW<C?\9XOc/;5.d[+@9(O[#U[
QQ_/=CPgLQ@RVg08e1Y?O3=^8.IU2D/G.FF(F-N+O&VIX_82a.:AWS&.A_VTSWH<
M05.bG:OZM:f-LMNNWeZ57cW?KLM4;VFQOMF9:?a/bO6:^X;F8/9W33ZQF\5S:W4
\A-9HB.+\AP/-0E4@2gYT>(ZK=_V4S34=X&CC()e@L>+KFL6FD050&D9FRL:G&G&
<TB1cM;YaY[-(<1QRUCL><<9+\<R17.I9GY>],g)@g>/,7#W<RIB\RAML5T3WLWD
72-=BIG;RM6a06\\B7RBPL]QE(U#^/?/IQFEU:_#TdAN#H)Q/8(WIR2X4FFMcTI1
6;X6b034P.9(P<2g=GBT\(IO>YH?CIKX0KHCMP/0\@L2RJ.O54PEL)-TCS>Z7+K5
WdGL;,UEDN@2_L4?b3IEVQ:-dMXd>[&H1aAgg1d+0T^9@LSHLOM\ZXU(K;F;K:-0
2_\VQSV33;0L&C;BdJfCce#_[fXV1NL0EIcUM)K^deA]^1Z^-[+82+SQ#Afe8WWa
ZZcR?<0aE[Y.,UP64#DRSE:ZCSg7;)TX?c)a9RJAYDH#5;R>K8FcWVeJH]6+>B7_
Ne[>.F(J(24]N(JJ0U_G69[0bLaMBeMB&9W<X)-..64ZF106#L4=M=VaNK2P;;D>
ERCF#KFN4/P\AXE6H3/gJV>_P2UfOTO:EVQW<YAFeZR_f#><Dc2>QTAaAQDEB@XS
ECP0bO[V2F:EeZ3XW_9/,]-YR-:\O;,5^E1CLR9L(]F\/TM)e\H9WM_WU(Y\;M-S
GSO)/T+Z>1MWU>C1F_#YWA#3g\:]c&E,\U[b\dQ496;C9#bI04;]BCI\Rbgg/D#8
/+YC?2\07c5SU1?cXY>7Qe,;>I7>GdgO^@>ZTIgAa81M<F8:C\?A@F2OF#XFGSKg
R-:3>7&Rb\b-N9DMLF6KPS#O>-4)R78J\&TX,#c<.=:.WN7\:&5@KGM7_bF7Y17f
YRKg/#1C0d8O41Y<M54[SA8QSeKeD=F^?S+J>cDG>,:(PRWRc70MU@@RA?ZC:efI
P-I(O6&[7[2a_>J97^&IJ862GEFP>aV]eD0FE1R,/eS#)\6YLVD-E0NT,Z3J5bXG
Q)B/7OMB@,RR8V0Xe3,/gd^9SBMEV0T.<P_A2KNB0&3#OTDf).P6f,D-Mb>XLeCO
L8+2SQK8<XOgPA/B:2&0]U-;c:\RQc1?IWSE>YPUCcD)L9@7+:[>)I1^>(5K\g;#
Qb\;Q8]Z?d3N/ND79FJ:TX/dKQ8NC&P_a2V2OL5O;P>\QA0H<>=E1=-97M0<X?/V
_f1G/B#SG5S;8e>4Va\JWM2-fIZ;]8PMS5.X3:T:^TR.<f>a:K^6/,Ha6Z9GeT:H
e4YNWJ/_;A(UB)<Z[QCOPY;/G01d#H&O.f\^Sf<Gb@KIFTHU<Mf4WcJLM@27C9^)
Z)fEQ&8I68\8EeS,UE<9DEM&.c?K7_YT4W,#DQ[+B43SPT9e#e_?2LC+QK;>cc,N
fCB?+W^=46=.X2O@I,W4ZDX=c+J^1Q=:<=@9K&,W_\TBV935S9F;E48bNQ([Z9+g
UMIfAVR;E?gM^Y83RB(Qg?ML:::J8;5+I;-f\B&_+IQ=2&g)7]W@A;=ZZ9)&O-TW
V6>N+APH>++(f2JIgVafcNJJU@(&+K(0Z9L_V(#_3]XJCW/[PCc]U<g<UW;?^>R+
S8.WSBfI3.<dHSG_I-Wb:1EJN20CB89JcTYM))@@dM/WEE4OZS)=?=:X>(OPSd2.
fM0fba9K.a@D>3WT:7(7+4+CWKcXM=P:P,gUG.Bfg/;A7FAQ>,0/TaR\QV<@DOQT
=21UG.+P5&>OSB<89a37.^1ccT24&+[PbVKK\7.Y)99PY1#BNC(A>2YdC];D<VcJ
\g3]T;[aeeL:+GHBN>9ZXEEe[XYWP90<>R=?&W2^b<.O5.eI2a.FU-0gM>b0P]OB
cGJWYg4X#Y7V3LB8,VEAE,\K6-g<Z4=YTd5W]2<5TN2XgQZ-QZ.JcaX6_b=KW.g@
LWb)V,Bc:B=AH=PDd70.2Aa4R(0eWgWO@_4CNAER<#>Z25e8:KXI3)4ALF7Qe>9^
^db1f2BWNTdCL:PeUO>AMfD.WDeg:_CE]?Ua3W^A/bVf9)1+?4V8]Kd],#?,P&PL
:b6Q@\YI]\NRQ2P(2K#?IdAS9e\.0Ra5F4=6-[b=0I3,:541MS4W0?4B_A\c]#QQ
-LO</1HU8(Q<E0XX9I?8dKC79?:VZ;GWdF&:(00.Y,:V.fe\)VCf0WA__fOS9IMQ
V-YS-A6(ZW9eRHV.\bV&I(:^O<,c,H[U4C/bD+e#6LdXZd:b-TZH63))<>ZUS3RA
<.Q@##(CH>dXMA3HJH7.^J-d=]/@]3LDDRb4QR,16KXUP,;QRGe>33_X+MIZEfXg
3V]+_;#;+^(K([G[7DLg\CCg40N=ER@?^I:R97MZWI][6cGc_d1NG@J#>Yb:BfW4
Uc\04HMggX^)J:]/G:f)R(CGH8(KXVJ./1K+QFE[9[BN&M5GH9,LYMfVec:=6_.<
\(-SfEc5HKgNT3[77I7KO>(@Y0c1K2LcLSOBMcL-aWXa&ST=W7/#=VGEZU?/Ac6Z
I?3e_D:1P#cAI(4_NLX8?4?_F,2f]V7))e)5GV35C^TQC[/8g8/b0O\b;1EIVd#R
F/IC38JYf:+D7Kf_8?4eNUf7R.^/M?.\VYLX^E8GEe&8bNdb9?.eOXCH(#[5PANG
(7W_QN(08ND59]OQ+?^QAE2Y6_NNBC/[GZ5=fH75IW:6-Q0T,.UB<EMdC2ZH+>a^
=;<^08cQO6_]<-+JY@@O;e6^G>0;1WfRXJ,@J5)(3VYb(&HU;SK6M4,6(/LC2__\
:3,7T4:Bf2&^CF6ONeEL)f>D0KKBVYQeSU/X&5(][^2]RPDO34LdcT9?^PYb8gEf
8V4/QL0]Q-5O8?S:WH9+CO1d]f<1VN)&?U.H@\,V^T4N9]eD+E\TO4Vd^\:[HG9Z
FLb:01(g:-2;dZ,]X<OW50>6/OLX[bN5,VY3.2;W3KHJI:Q1QERQ5Y_8GT)DPW7S
PH+=a41FN<6A<@(@g#a[Y+GTY<Q6Sf4:)T#9e:SM0<U[YZ3@SQ\IL5+]1BPY#D^:
5UZ/;/bP]QYf[_a[I+[ZJ7B1]89;b8c]Z^YWYQO]Ae\TD,Lg]fQ;1Yf,9&::S,.,
8b@VX0f@@(,CM\UNU[:Hd;V>\)R=Y=06(;-2,F]DTfNFQ3BaRW5DUX@2baUECQ<^
fY>=OeF><0S+Wb@9g.4/F^AEY9BIJW:fJM])Re;gZ:\P)I-X6a@gWN?QJc.V(Ff_
=46?cO,[#BK@WeYYXI3f7D(/V6A51Q,?;:d#dC^S&\LJLBFg+M9&YKRPeJRDD4<O
@-5Q3EGTFg;X7E_ST19CM68+A8:#D_d=L30+fc9BP_\PSY\HU80d&Mc)=eK/BG<Q
8<BJH5b?@K3XBA_b0C4O9^C?Q&5b/E_cD^<?OSOQ=cb]^2&(:A;C2:4bG50X<#9T
P_dXY-ADgH)SITd0gG1S74Q&c3W&?61eWG<4K;0LGW/:\K5;S3+P6:L&b^M.N#)0
P?),Z\>HQ&^F^Sa4)K3R<&6f3G.2,]3:Y7I89T&44BY;[BV]cP;)?&=4b0JY\1eY
XS]\F2@:&-,\Z#GDX;GZ>4WK4(F@\@G\JJLY?TY\]O/_dQEVJ<<W5ZbbNB1)#^.Y
WV)I<6(CUD]g/O2eNSMJ-7+UJ54_L./a/LKHE^TU0:Z1F_5Eaa56g#]E=e[)aRL]
4.G<_R[G@&?S8e61/^Bg,DL^eS,K#FZJ@38I/:.3T&E3#BSU^,H]6MLQ?-fZ_O5e
KCa<)_N@46KD(#FFeEcTFYCCT/KC]bD)O+_\C;EFe2G_3QQ8?YG1C?^(^@O?A5L(
I+\^C:g6LBd8J;A<@bBL0N-fF8PYDS1;dbe9^6]4Z[B:KPUd]A(-K@4B)P2XT+.:
Xg[LHE3TLUHC=^J#QUP=Z1fKXD\Ff6K1I\LB;0,Q#0#<Q:^HEc#M6/D4,_NI#P^<
4&)+]0)5bBb,913OHTec:/2@?YX\>3D<,7<JA4cE_3+H5,4eDU#TcDgfYR4<B]QX
NU5ZOUXLAR,KDHI.egWVG#H2D(;WV?)b8,DXN,/)eEZ#:^.KN#?2^5PNXgX;Le4T
BV.>Y:<6_)c#JHFEH6/X@6b)OK2U=3_T7BIV:<3()gNf2da3];5[3PdNe@UZC5@1
1_+P\2eY/3U88a#GIQ3S.B^.JP/SHTE\3cC;>-ZYdT23/A<G39PIV/CX766F6@PQ
#S^P[3;2YJJ/BMI-?K;4V<d95&=R65aK=WUf>&WW^(LdFZ/;3)^G+C/#I_:2=D]c
D.g\PD<(8\9FMG[V(@\?-_,d4f+6KbTQL>8OC2D4>gM\<#+?/15[=>&47OZ;6CGd
RP)]8#T-+S0<WF(R,Rd8:A-DgO+MUX_cKCXC8YSQ]H1f.C>SZXPd5SeQ6)T0H/97
dg&2>KdRdO+00JOAW<KF[.S5g9TSc](ZU/f9T1<D5,HUDE494#eT2J.HFf/B+0/M
BM@D:3?7&E4<S,78NFeVPJ-JcR/J>\N7US.6Y=QV&gQaT[H\2D.F-?)[I_0EZ(YX
XQb+4f)dd-@Z2J>8HaV3_<IKEO[VGdd=;08aMgCQJNYJT6^aYM&?BL#KO?I@([-Y
7Kbf-@D[X_BDML2,0d)K,\?7\&A3D5L(6\(V^9S9#f8G#Y?3S?&X;6R8Cg^B@5M1
#&S4O&32J&PbM>GV^)5?2_0#EH(JQaC,@a5ZGM?J@K@0F:eJgE]fKfTIQ^b3>4>:
Z@&9F//0MbCfT6JT5EDdJB0/^,8fQBUPZa5[&@b7B_g,K<M+>T)(4bHCYB_B\[T-
@^T0H.4g^c-<F;9ZDKWeeDeQP4L>;:7/H/b53,8(1\3]+VWI_e(eD+(+2VH.M.@Q
O/X7P,^a:?=5I(_-a>HIL7+H)0Q\D?\YB;;/J,C>NM_4T2YEBS;BJY-81_O,A]3+
TS@#CfWX8>QFGY);^cb9WY(PZ+E4MBUJU@1;FML539.B3N1:6<2FF#[U.YZ+DP#Z
S@1HP:;c4]8YbB6@fbb?CRL,?XfWRNge@XW;R(EBQE&H_.J/(4<LJ;^DaS7a^/;Q
CF#-W86f_V:.F/f54FLS[&N&+5(A[,Q_Z?^#YEEAQ8D9;U0f1;6^:C9DbPX,J#gY
;W+&85:a.W3dG1c8bH#dc)S1_BSY[aE0d._?5^VUV+2?g+)Q=Hb?HR-MMc1J,F0,
d/5).@d?D;^1J2Te#R[J];,?2F.;X-JO?I7;Tb\H/\.H.7d0\18KRICg4F<UVC2+
ZARIIMFV/JTR<L?6@#@EE@cSPIeHT6IT:AOMMH2^W>4^LH/I4<XE<a?[gI@,e7HG
_BCeHYPSI].9c94ZYLbIAFC8_Z7=.MRIXC5U^-ZgY(dHP8@)LB+a>W@Qg;<=Z[6g
cWU9?KT1Dd0GdTX1]-7]UQN/W-4;V6LLgTY?Q&4?UCSH,B7g:(/X]TS<_Q>aD0\K
c4+B_YY&9GXcBb)eS(NOXGGcaTX&EH3.,S.GX01c(1YTLN#I=5>96NZY4Z;C7U>Z
f(>F+>?+IN\O4YI@F#NC[V2<1-ZSU,7+O^&62ca(UGYa&bKJ#4BO?:8H6Q/MAPVC
e>aP6#NFR#6T=U:H2P_VW(V\]\c<gSMIVD7A9;?WAH_W@L-P]\9FD^WUF96OUE0b
K6)X\7AYZ^##9.+(P&W0S,M/PO]Y3TK=d4cJUT&bf[VJR#.&_YX8?SQXY47&K/60
Z15Q,PGQF^JQ&4>JQ)@fF5PdW5Cb2F8cLf[J2Dc=WYX<a6NJKGWe98.#=.U5>fE5
5S>O^JL<9S\,<P27@G<9O]:E?)ENJ56.47=cWN^O,3Bd3<<;eDMb.bJZ#H/OSKJF
<GF3&L_&g[@MA.Y#9I3)agB;[c_#\#g&PAW/DJ9/RL\Sb3?VXb:3G7OL7FHd3];?
@I8G:-,/LR#]bD>>K0TPgfX,d<U8IeWZBWXDdP-?313aeA@.4JM55.,S;Kb6f?2b
.cX8#_0=^,,]\GD:>f07)Y^=Me7EQ.+YP<FPWVcbY8B-2\OK6R?1+F&GYP1T-NUA
N2d3IbUPe:CM7DBE@TLO\1c3aA:N^^M]-bD#+Z4N.7bb,_@Yd(.IQI0UaCZ0<)+g
6NBIYQ;fXG;b-+YDgCbQ<R5Qg,P7@:QZVcPMSY+6U^[]e7agL4Wb#@cN\6>G-ALA
eKU59_;B_&T\_?b0(IgZ6-N/c[b&Y0)S@+WgSf?8#47a&C7I<:&9GD3IO./&)GfK
((V#N54f:RJPGJ1LC2/:>eU.U,1JA]3R(R\)(Y5C[WEHg/>V^d7RK,LI^aUUWB7X
C-S+,;ZbgcRC>-B<ZSJX1U[GH2.^)5)MH1U\2JM<PMK9C2eCV2M]IVB3cN,Je>(G
cS&V_(K^NAZXD#GY&Q-<C+/M0_Z;gIO?6eL7-1fZg&CG1]MQUBNBDJ:44)F.B4SY
0(UTW.YL7aNIY,GO&RXGaaN^T)gJ(#SZH@Hc35WV+caXJSSg8eOPbWeEL&7d>gT&
9I[/+-H(V8;8)8I^cMQZQ-O?[3M-@#=^GJ^OEQDeKPU5TQ0O</([4a?+NL@LPb&c
WgMWDTADFPB.0H4:N5RG/&DU;IW2-70?D]=dVZ<8Kc;^IQH8gWT#LgF#BJTLRE//
-CAK6#2>TGQ5Nf&7e@14G.2WI&a7+WDeC98F?11I+5Z+D(2D,6Y=FLMfLDGGFCT@
aUZABH[)dO,2f-I-cIVX7TZ4D9#[K_3WHK<J/b,056+)U7DZ\Kb\[X^@#gRJB_Z9
@cHS3F5?^L8@UFT93eGV>Xa;4bS-f@f#3_>TeXT8Q)U)S-?R)_Zc_.24K=OE.Og\
7THRE?Y>K=GY7_PKCL:.G:[Q2N:EP+[UKV3T9IH.0KQC-f-fX/5]+gEY01N;M4Yd
+4=0,(KU4>9/e+2^\Ec>?PcF-acD=G<L#^(OJc+V_PgRe7H]e\AUY:MRA2G<RVT&
Z8?G/O0^CTGDO^X-d2[DV:&,NAC8BNGfPecC<X.O\D8a[G:O<#C=4VcS=[DMg2bK
6-:2>-TBS)?/:1F&MF&c/D;.S/Z/;I)f866O<?^+)Z5C-985HVd&.-?KU1A6b7SE
EbE#MW(4VC2)H^ERdUZ4e4Ud0+9fJFS_;OHc+;#CbA4e?UX?=?@>4@E7.G/:dCH+
cBa1TQB.ST2:=[=L44dS;M<6]E?8\B5C=CEY-92g]JRY]6e)J/R6cK)\OR0a_UBE
de(<N>W#/>18Va4ZTC@WTYL&/2KE,BNECQ.T_bGC#<5FL)2J-\X.GCVNX/A,K3ST
BBB8N+LgGK/P.QB/aU?S++XB+.5aYd?PO[#\TI&ba]G[=ed3+\?=R0&M&_\B[H(8
3_K</&c?K^TXgbcdcU5B0/fB&:bV8CJL&H1e5F69#:[FRU/49XbEN,9A<W?G:U_^
K5@<YWN,1F9g8(F;N03(?9L<-&4_C@;[(4,2GV\.5_.Nd..5[XI?ADZASLC-1,34
7.@G[aP3P8KQA\[D.Q>ZH8<Z?;CVDCYa\X\NF>QMgIc_C^Ba.<+@NM:-?2eB5&24
F3@7-B:DF+HJ.H>.@c_PeLPg5^ZB3Cg1A6UK9FR340BW\bRF(1+5854F,XK1Edf]
+E.)T5-;3TOU8.]9-[O6&N9#FXOc/KKZ9$
`endprotected
endmodule
