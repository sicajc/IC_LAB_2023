//############################################################################
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//   (C) Copyright Laboratory System Integration and Silicon Implementation
//   All Right Reserved
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   2023 ICLAB Fall Course
//   Lab03      : BRIDGE
//   Author     : Ting-Yu Chang
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   File Name   : pseudo_SD.v
//   Module Name : pseudo_SD
//   Release version : v1.0 (Release Date: Sep-2023)
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//############################################################################

module pseudo_SD (
           clk,
           MOSI,
           MISO
       );

input clk;
input MOSI;
output reg MISO;

`protected
>4:62NcIH>Ub^W<f,RCG#0_<YY&MR?#f\c/>:4M9fOM_INbS-]774)?)I:&CLX1;
4A2_d4OACDCD1RS;9Z4MEEIB.8)FTFAT]PO^JedD._E>U_6A<F\X_5G_\=;X8NR-
B_c1FDfH[JTZ/_9AgTE9^H(KFUfOOX3<YL5b21)7]WPNKMdYccbc>C>7:(3B9:dL
AK:cZ;-0d4EKZ29+QL[eZCgC/IRLM1ZWEJe8]FN,3W<OC=9>f.T78JRFX:5ZEP)J
>KLD]561Z7#3Ee<R4T?<7@YVLNTUa9/,_D)3B1F.959Z[JcgICSWdDR#-9,?RUG_
d2&Jc2V.I(6=R9].fO.<KB-N9g@L[2&T/6-V&;[A(><--#H#_Z>W(eA=XI2IT^D<
_+0\Sa(]eUV&0ZU?LdHG9+V4P166G&\TOG8)&Q41a2]d<[4Ja10UW4#,4FOc+W24
^_ZVX^DS1PfcW1H7V,aCPV@G-I12HZWZB=W[&#A1CbQ[DH3]]2S0+K:0,bV#Y8\W
MQBS5QM]&d=?_[0NP#P(M>GMW:X&R6Z9BJV<K5VD+-E(aE>2/=J3./MI&YP-09PC
6MD\HLSH?HIT>\ZB-&+XP+J8>R,4SC&FYI)10+T\Z2=/<eNFQCJN3[R\3J=Z+(a0
e=^.;60L^Xg7Q0ZgO107S\TICR/#^8/\9NAJb.S].P]^XC(<D->R?--B@4YQSe.&
5I+MeS\,a8?B__\MI&;U:,JgC[QB1LMN=NP^43;f9K/ab>&G-YM&<6F[QBS@MB)\
9DCIV#L:Hde,:9fb:LH_C@N+G63;K)8/T464WfA^BT@>9#Je7T=<14M\,A+-B3#B
8][e?JU1_Y].<15^=/Uc8\8Z1eP,A30f.?LI5dBU^)@OFAVR\:g#D/)fA:E>9^I4
/JXdW@<>2@JG6&e3/0AH>S&gGOOcH-He48b>6ca/?Jg4G&J2=Ud./G2D-\c)NI&^
6J?>3(M@)QEW@^6@AWUH8==]S(-]?08b<\0J4/aBg@#fG<M#RV0G1#PggOPb0HX]
cg.&(N/fH,YYU&a5.CKS(@GBDIXCKgKON?I9HGb]0.6?1^2.c]29b&X08cWLL8MV
.F<PO=cN-1S#O8XQ>0]=3BGBPHeX-Y>IK_Da.a_R4;b_/I;39EJaFF[06+O06eg>
85-M)W)9#-G&=fDOA5S2c1RD<7W5N:b.6U(;fIa(&Z:PO]bU\CK5^dI3Q&?B9[\^
IHWdMZCTd@HBbQJH@X;3Y:D;Uc0)JGDg7RgNA:\I=gVbXd_eZR@aK<56NZAU?E+&
EN(3dQ74_\GZ&\5E+-4N-.JQ,NF4?>bH3=7c=Q;O(?.1I5GW_0f1F&geGU9,14)Q
>>VMRUU/NYDC;NR^,KI65K<AE(NR1J=9cSDO_G6Kg-N_WB5eVZ_;C=aN^BS?[b)5
]^\fG]&STH\Y=<2>H4,_U++N2QOP=(/eDMP]Y7-WYT;K6M=OB/@RE/<B,W-Mf5&?
W@CF:-9C0=@LK1ePO/<G-O7O#.ZRJO_R=.V0-&+E#04/Sg-C__eG)M@?O=b9PVB)
@\L;gba0<@^eL(K2X0=Af]=;3>)9g[\7:(5=:WDO5NbD9aLc>&(;gY+I?&f5.Vb&
GBaRd^]+cOfC[.agbLfG+AcbFK#0-X_E2EA7&>+I&L04RAUD(:RB.3AS0aIPH3&(
?]J72V&6#?/bQ[D:8fZ5dgNI62T8^P(Ab\3,Eb<(>QKC-5W\#FT/fOd\_XG@D=P6
e<<Y\<>cKM]d>2cIN&2PMYJgWH0UJ9O-QQED8e5@L)<dQ9P[4(gG/]3@)6.8]9BJ
<6c-3C11:1O(YAI=\1.fY+QP>L)7Bca#Qc3;\^9/+=b]X97gI3OR@E,M#:;UK)RQ
7#\2aTG)Z_TY\TJ>UHeO\+]Y72CISVK)9F51Y0)\5OO4c0eg0=cSVT4(U#<&^6Nc
E2Y]RQ9Wef&U>cH642QN(GSg(]J50C_AJ.U9D-LPS]^BMC03W(^f-IJ&PFC09MF9
>7Z(c^^=3GbGcBL-g+R#)ET^c:CHJSFM(8bJ>2G1+aC1&gRD8QaQ:P2Y6N@cUGTd
Y29L\/cD>U9]FbCBbZ&G/RP@4:Y.DMIJ5]aTPWgSM]Oa\9Q3W69I(dIec@Z3F>AB
gD-].S4M/Be2:;6+F7#K^\O.0Aa@cgfM/V5>?W8N/1_+@PANFJC;[-0C#;6NZIHM
0O&a@?K7fO;)5/Y/;dOA?bCSF(@SCR0]@_1W@PG\(3#Fc][XX(RTK22V7)#OR18<
DebI0Ga@b[JV2(A.H6WebEMOGO/>^\.)<Gg(,09fg62.BDg7)Mb->d+Le,0Be[VT
;IgZB9W/D(dQ^a2dV7(RgJ0.?;2M9<cQ9N[YBG,]J5^)(99Y;/g1f63Z/)P^aMMU
J1d;Y.A1PBHHd<0[bC-DTT)YB,ga[?=#0XeGePMIS3cX-U_QLe&ABf@+UUQOI37V
&FLRK_EeF:G?D.ZI:/U+N_]W,CGOHGcO&42&d#]H-.77L,cC[Me-(J/(=IGd/A-/
DaLIJB=<[C@AQR+MT=dYQBLI0A<+ML[0FTK(>W<-TY;Uf0\1/#9NgZT(ZfPW-_Pe
E@5J3/#C<C;gDR;(.A+6SET:]\gH(4\5^]a\;+2JQ(35^@)KMGK0TP(YW)<ba)JW
O[CP45,+=CT@EAWUbJ\9V:J<9GXJd1BgZMOG7Nbc0C<b-d[ecUfJ06>T_X]D4TcS
E0.[7Ode>C1c?AM7NX-(G]>TF+.C\&W?dS]2FE>X<7._YSFOc?#[Xd+Z73\&,LZ6
dX(GDHYP9ZQ=4DD^J@_a1I5/[3>EVB\Rd9H0[ZD#d9-T6H5DH7GdJecaCB:5^.9D
3;&+:Y4)Q)?8.&3;WM.(V-42+AP;;@eXF&<,b;2P)_BEf5-H//Se88G>;eM^]#;)
J@9?3a@4S]J1?\KMJA[J;gc,eS=M_Aa2?BeT5TPTZ3<M+4;RA2L7N_QQEDASe9c1
K+cZf3JCEdU_RL^FW<0OFKDG6LCTO7:X98PG[K__9SYY[XY?M7b\X:VTcc+NHE5N
Nc]N>;a7a6(\>H2>4Q.JREMH5b#_)eebQAI,?N:b0U+V;1CC)]C,Z3DXPe=R1V:^
G#D@^0DKY9E35Z91^L^^^Lc)&367fK@+SJ_,X<;3c786]YU1dX(MK6WGL,J>=[?3
8g3JI2S@T<0ebZ3FMHD/Q^g)BRIH8@F-AgD=LU_2M?3&=];fVK=#Tf_?^MG]^bTV
T:9V]-Gb5eER,H,E,^<:Na4+Y8f;Md22NRa[.(6_W0GF+BNSP@dc^G9LFQV4]3g4
PMBLC:,A#L89,T8\a[5G(W4:e_GC^HbIVB(HW&]B88P35f-<?W@?>F\-@R;BZ]J3
&7aJfWAf]02+:e/M>)XGL?b#gT>AYMN9U=JTJ7;f87W?CZO+WM2_;UI,a7bL8dWd
,]FdC+Y3S-(Q[6F#E)@fOg:=0.M/DSGWLEb])JG;b..9[4,[\#A-5/<LXZU:S<O9
HC9/CQd0@\&DI8E43LRd=SS)bPX-2EfMa6XC)L91&3K;/(S2g/S?/TA^(D:;.#3b
3KMN>_CAC9XF5-J7GM^aX\PIf^b74XH;#JQa+/&2eO8Q]3c^Z)=0g>/aR,+Ee&W0
bJJ344^eaJ2)2D&/Hf?Xf2,W;Z930KI74=@V+_/U&PgP7K<LaAJ6bE2@G@#(RXAS
a3K3155,dA;B4cE^+bIE]D(D4M;gLa9a4]Z@ELcB8(3:(-(OFJ=DB(\(Hf45L@3U
PP#/V>9UM70-;KKWCJU/[Q@U;b?>UIfT>6N\:F&)=\;T/:\L23F7Hb#9+Jg=\aIW
+OLD&fcDJFAO#e/,&KJ=BFR=+.4YP#FDW=3]c?N7c,P,4VcY2[&]:cS/,B#C:<Yc
O\-,:2HZ3eA#fW,O0+=3\^P2XcD[+e;]2UBa)M#5P2\ZdI7.9aT(Q1)K(YJ4_Q?S
L1=+\1[)@(0-cEd\G[_3gOV1<cP4YFd=dCS/-3)<a6GeMS]7bC6Ca:>L09/.R^cT
,@Q/0,2Hf)V=IY:V?/_HH/>7W<R)]8KS4W/DUO<Qg)U#[+7E71:#BTZ/H+H65RG@
0SX/R[LZ&8>6B]K\:+]&HJ5\a>N_L+ED5cbJ,SY<c#eKOfS?ES@MVUd-M9?)/8OW
Vc0P5)[93.[=-U0VCgR]UUI;:V^C(?7]_GG2A8QM_,=WC&=-)6\<]JAO?J<R+U\;
]ENMA&;\4E]Nce=/)P>>>?L_+?D^[VQ,aXdJC0W^3eGT/J>g>+Y7?:_DTL[LMH;B
S<ae7FM\:8H:8GEM]?gcM:O(aK-2W.A6X8KV3IZ.GL8)(H.g?YY4:E_V#FTaZ:(d
-)IWObSCT);MM4LS:>N>DaU<<9IVd3K<aQ6F/^DQTgWC&GJTOeG)eYK0XH):P.T&
V>;<1JNDQY+^bF[GR1@fY/LgD_d>(+4QO(K,;QN-O^_H7&3>\SAGH3\60>?)XS=J
>,/c+FWW9Va8YB.,ZU&-(JCU<8&c,W,_[_Y^Q7ZGdcU.7QQ:L86NgXX;/DEQH9G[
EGYQX+8]\?)?6_35;UgUX6A)L=/>cZd_?8c/W+XMLUdN@1B^BX(4X\CT1a^2dIR<
1G_JLK&#)/5]3?OY,>YD[^K;F-:X4\c5-cJG]#KFWVF_@3FAGSQWO;KI1K)KD5]1
EN@M3;C1\NIOZ_](FSIT6(eYMBH7\c6[GQAC9>g<ZSW_#9T_)QQeN(dME[S63_DS
Q?B^\Y?2^)&E4+N10eQ_4L[5:Y^eNaC?f)9fg7cR2,0^#U<>AN.dBM\G#TCa](6=
Z+/@TE+P92TA;3a1bdL0Z/S1V5Q1gC)E#&0Z=_TO:N(0E@4K7?@J^]8@bXPL,A)^
Y49/3bRC+Y1BdbOG+,H+R)6^1\;BVRO)Nc2-gT,5D+\Qc3cH[7bNR\4X>R;AEG2X
C<:EH+0GSPE10>6EP?F/TU3V3.6c<M(dZ.PgVLPW#^aW>HZ)7\W?+#fE14IU^WE7
79U+M+6FR::bb,>>P,_(S;gSQ+KYK995Xb#b(/.aQR_DU//[:04@8eDM+d>:O;=g
G1RP,.8GZdTSF<\IEXUe>M+dX71.I1gK#((W@3,GR/B\BCB\TKGD#H/1<0D]<aAQ
O<)I+bY_>V6^-E,V>b<Y_#LZ:\eG,;4#SC3EWcXBWJHW13G=IN)Q<9?TGMTT>fBc
5eKdbcZ(Pc0[fO3]#gRV^?LU6WJb+A-[^)gf;MJc312@a_/#=O<e4f.TF^R:<9I0
KF\<PFVLcA.[Z6RM;](A>c]>aV7^UFLL_WfK)#&+=:eRUIFgVJ@&002G>[?5d-L^
-#g=d<=[<09e<WXBH6:aTKdV]C-GCLb7NEb(6H[J28PcX>BZN^2];G\X9f[>bE)O
+@B4c&eA[;5F5=/WXB=g\@H]M&Z-(IGVCUW0WdZ5K3a4e;(\__A7G6XfHU;<4GX]
#_@2;T5J/2f7CKf-L]A29ED\bRgXG++HNSHefDaWb#8:aYIBAMRBLEE@BI2TA5N3
,IaHc:de0M^P@SG9@(1+d9E=&F5L0W3Y0&GYNP[^81-0A]F;)]W.O>VUVJO+>0C_
3b7VgQHH3^If]CaU?I\@C2>2JIcX]-NKf@N:5.7-_XgAZX)g>ANFRPS\[CY>f+Pg
_F^g4=fbfMN#:=Z><UE:WR0a5E7I]M,]WXb7FTQ#PG1&6USCcD+>9INGI)RQ9<M?
0JQMD[JcZR5#/#7eL^M1:3dM8<aHO&NO:_/ZX5HMJKV@]e+J0P<5Q2+cg?T2H#eb
I\W]MV:K4MG5/:;d>/aREKZK/XYDAC>4?3bH/6@eTTR@\-]N+)#S7BaL]L<S^B]1
.J/-VE0H-X>]M,MD5-F7>I/\W^G9&:&YHeQ/[=#ddLR^FTTHg0#46OY7g<4&?\P^
)0Z<=RL^VFf69W6NMe2Sa3PX_GN>-[F\X=SN0Y_SIT#d[+&-,Od.Wf4S^d5B[fcL
g7g]d82AD\6[-3YAA3PL3BcO,S;.MY)f[X2(;ZV&f&[9DUZ?8D-XdTK<b++I+@6Y
>g,LB>2B8EaI?=W9Z2,J\4T4NOV331CV)([JcMWcR1URC:3a.OF--3@,Z-?#O5.g
c(EgTZ_A/_&fEFU+^S+dP]B.N0+)0.#1QEeY.IS(a+c0/bO=CE\f@WR9a.1U/QJN
?L7(.;;_Hf6c=3/V@&cRXeNIW0&3F0U#E:@VNVR1?#/=Sf\&E()JPV;FWM2(0,Bf
RC+3RK1Y1:(^W:4/>@;2aYQ[6A2/53LQEW^ASQ1[Y,g[>b+.?/2a+5^20<G9N,K>
B:d+DET+KU_c(f;QSVN?e=A)LHV#3FM0+@TC+T,4GTZO<F_&U2RCY21#7R2)FGPB
]_g@NX]-:1-<]\(:43E.4Sb7H[R71HgW[gGEYeZPZ(:KC4TeYf(a:33RA(&H:BKG
^[\a/daD_DJS\]-C3^PA1c4XO^Re-3000)Q.Y<7B=?Z?JXO94X].A(VT@Y73Z#^T
D6#Z:-H.3N:OD0D5J7NMFWIfa(I7MXSX[fQH4a8RaC.Z:7[#C282;Hd6=W+UFR9&
]WXP6;IB73.bC(Q&26UZO)BfT,^2_]G6(&)R)TK9R>CN;;N-PQ1=a7^,6L9#OSJ5
bEZ09N?XaXdLAYgb\)]AH,P<57YFbB@P5]6dFI3K1EA9/(fdCX(72U5L,e\)X\Z7
KGeO+bR]^A#A)L=J@DBHGBDHfO0H#00+_=3I_1CRWd]1(V-:N,0>S\HM[F0c<WX6
e.4,1=F)BJB&1IbA_SX+G+34/(dS1Jf,]6@a/G,/<8D7>K,?[72.d:b/;1IWG/H\
1&9Y4OKP(Q(T:AQW,1QN4NLFT/ZcbGeV3[)5/8;a?=;ID?;=2?67\0VD-?cP+M;:
P/B-C[;eA+]:4Z?&I]UFCV;[1HMV+?4)<F=1g99gTL\;bW2.V,#H?cREF0U;=2GJ
V-OTCYc8/^V6e]NgMJ\1&&AVa(g_(CJa.d8,EC-T=(9/Z16EHR-Z-Fd5e&eG7?8;
M:F0?+Q</XU,YE+I[HO[+D-EIg[MFH.]R8+70=G1#Y5Ta<bg52=+P[OSCb#E,cC=
:K>J55Z:=O.;0f_,/Y3RABB:2&\+G]/^]C<<P]T_UYg0&3cXbIGeXQE;2/Ne=Ya?
#CR4]4UY=?&c=8-LC_8)(IQ<9C9[HX^eA&aT,.Df^B(PC,0JE80_A[3e)E@LKdAd
aGIT/]/DBT&d:2S7\N5bM2B+GJW<f3WFcfO4PgbTHTQS7I1WNf8c]Q_/UbYBcg[C
23@X9/1fY1gJ+F+2FW[<,C[&5Ua-b3P)K7FG[WGP8-ET0<2AR;>K5ZRD[Y2_[MRP
-(L#dQT(^:G#QdbggF5SGW@==cRb413I?H-R?()T5Z;eL3KMIdT5N21CO@Od8>_#
JfG-0WFJ?.P^WO+DSA,IGN(W1H;^G/Q_TH<[C[OW3CU4M.DIg\Kc>0RO0KTFVSGX
&)&57-Va6(@F#+J?Fe&e32HT+KNHcGN\eWJZ/9#ZCJU[(&4K7TTefY-CA;F&A=PC
6)I:(A9]G,g:+PN/#75]Lf11<eZ[d3&KFd,4K]E9_aQY^A<.LD>F.<;;0(_FNT+B
=#+6aPEJR&bTKf/(=>B59/S/C9UQ(4)\[cM=&:e^2XUGAL4&PYC7=<,aX9E.Q2O;
g;#V5gA&3cY+4gIN=Ce:F11Pb8Z26V^GFBcL3(#YCHU=[<g?<IXBW57=-39Sfg\c
6\O_W_K8POTIM?2>?^H&+#,Zc;A+T=<:;1gW>S2de9Yb3LAX,N3QS^V)GNFA5a5e
7:S2CG2^622T213MM[42BbEW1X,\-2CM#.2&/5PO:Yf\b2,BH^G4;F7O0FSJ4:+f
a6OH/>K@QaR<?gEQT&9<,M69;J&-EgB#e:KbEZ-RC6D>abX1X<[PD0LI.gcNg#4_
OK<I+\]CQVSJ@[:1-g;gXL4.^8CS0-R72OL?WLF:+=&LdHMZO1]aDDeX)=8d1f=<
VT\;fDK+Te&S^Ad;>_?QHC>;X.C+Kg87CJa_Sg<1U7&Se=_d9BdJ]D>bXT4/\GM/
U.=]BBZ6bEa74d/AI+5-d0PUKD+SG[U6dMEN6F\\:.XVI[;9KfcV?PJ7XSNde,AQ
d)=]D3KDYQ3]fRMF&H-&VR<BMWSE)?Q(=Q3+e8H30IB:H7;&W?<0J_:,6AS44c80
#=^]?FeS8DDc,1K.8F6H75.KU3aQ8.#aD.WZXW,N8\)PX<Z_b8G4N@c#^Td@2S-C
AGYB]\65<D3@GY6HXO/WPR,]B80N)HZBV.A#DI7DgHc5YPPHDg/CR2,84CDSRLY1
V])NF@PH:?W#M^3]]K&N@ZPN,M>>PP9IZV:0B:R(Gga&?=(B8(+QRFH7)Qe7ME#1
1a/bb+IO>O,8AQVJY(R5^Hf3)7;IfHFD6:3VJJ@^7CL8-6:UA,3R&3;I]D<TdAA8
JV-=gN#YeG@c]&P/.3NbZ;Lc9PfK6.Y7(U85-<LEdKKO_?CMe2&5N_BeMK,bJ^9C
)41]XBcdU(5-:\^BO^b@<;ZC/e)BLLCV]E;dJBJ;SWf>S<WG#,cd]AYW@bfSUZ6-
ENXaQJFBR-VM]f@((\Kb==;]<cV,4Ha=,+SX=b@WUFIIXO:^d[:R+#24&aVP..0F
TWdE4@=;O_-7MCO+FEfU#CT6Xb+Z+>RN,/WU0S_<&c.e8)MJ9?XAMEcT@AZ1_IR;
>@d6?f_/_gc[bT^],GV0^K1CB.e)IJLB?bCbM0V(UOW^\T5JLOJ(S2Sa\D7#4+Y7
51G/#R+aS^U=\703c7c&5dcHY<DGA3#[#8e<,U(e9Kc[feAL#>G-07c6=UX1gS?A
T+E2Z]XL_;GJ_H2fP:\/(S^#VSHZQ(7aH^D;f+Dd:D4LZG[?gE8cUd#9e]]>7Z]P
-3J80PK4FR2dP26Pe#L4#N3/^(FZ(8c]JQ_JAWQAHDZV;Ne_H/YfWYAU5R&D>5H0
a8GVPU54UUR;Y[QSLY&YRM9HNJ9JMAD]S#1b3e?FXCdOgIRTKLTKW(^W4eE)ZQc#
Y,Eg/-,>UT1J>M9&1U4=R.HBF\,gG8466Q3S>eFSF3@(OQVABHc.O^\1fI+>^86U
4d&7O48:1a?-X;dW/_U5OG7eR\8KSa-I7fJEb^2_J^d.O-E;]29P2bdRaU[,UP#J
S+b+SECMGBU2PWG1FA38G8U29GUAMXQ0G/4e@dfPVH\5)=\gMX.MS+;9edY8H0FL
J8XDHXfg913#6g(#P.M&G87Sa9YN>@,gO0[g7RBL&UI6@PAST#ADJ/beJ8;)M?B:
Cb.X>cS=eKYH=OQ?Jf#<3&=TD(aZ2V0cR>I/(]75CV5,XGaeC]eXDGW7M-,/1P(:
0(VV<3XC0290[0G4Te]ReZMJPe\]3=@d2&caDRWC>e3_ASf219P;9&S;V#3.6bNY
]eUdV2@#c\;\U<S?-(Q+=TG?/_;?PCPQ?72QP0:b)0dCa1DF<U#:,<dXQCP\UX?@
d8be3)1_6aAWNafaJZ^M?E7.8-FOKR_J@I8+>OM=H5O;0)g@HU8V>[EN[W1a&WX_
/KVg\\R_Z^NdZ4X:Og-D=5[/:b+gZ,XY2BZ-C<BVJ#1H:d\AZL[ND:D[(e5+\Q_Q
[O.^)Z6\S2R^e/T8WG#T-=OPbGK)LB4O>R8;>594RT3B<^TK&CcD(5H6N(E<ZHLR
7e+09+^=La5\8,eeDS\<T1XNe97=,/IQQ=DC^0B#PdAg#b/BA.P?NMTV<?QB:8U1
1_)0@8]Pf7=4b6RaJ[8USb4MAe=YWOUS,71.If[V\K[LGDc]4=I3L[M5KBcA+HYb
Y^=>=B\V7YA<(:Q#0J/D[BEFJ=5dQ>6(2TIQ:<JJD_ga4I#&#/B=EV]:Xab><,I3
1R?EH@N90;3X<CV12DEVRV:g/G5>\=NNEG1?PN2R;I,fDFfOI6);Z[LUcNHb0>QI
@O_^6S3Jc=D@BL=P+FGdX0?<c-1IGGObNC\UbT=#V<b34CX+XGf825,R,SOMX5<e
NRUL2)abBZgF;A[)0P[5@gM;#eGFN8bN@26B&]aG67F=8bf)RRPA78XXWU=Z]Uc4
0U)9MDcfSJ,3PA3P0HLJeeTc:]fD^U+#[Uf]YLHH)]^^NEN[>SFB1C]3,K([D]-2
cI1[RMI)g(ZWGBedF6.Sg@90^@9MT/0NE3.G\UZ;ff_/DUH3/@L[W-5^gR&@KH.;
ZfULPB/34/4/;eWGd+NBJOcPc-<7W^(:6)<].FcW#MXFQM:31CNO.=a::RU+=-WL
0GWK<;4#bJN\.fL-]WNdHJAfX&2D1WA1TOEBZMB[2^/RMNHI@A[?9Wa8-NVD8:E^
H@d;?@fPI8IaNBN?<4N)SM.592g&Ib>^FRe?QSMR)+RBJFL5H.4/1M]=(1?Z_ec&
bBZecdKDg>0-U72+@TEg]YG(BHE#KR.C/&YL>.c[QR+Bee;^/_&R1/a7)d]05)Je
Fe=ce7=@<)BB]+AL[Lc[[f3eE](C9F7]-3=8U\@)D)-gb=cG#]&df?W&]9RA+7fb
@0J&S(e7&38H2Y::3VMcLZULO?N1G]N=_G1(0;P(H==6@D?C3WYT#<OS6cB9LEAH
O@T/1^SWEa3BY):YX8GK[)O;GCC2NMZ#W6KU8@a]Rc[=^2X9bN_d;c-72#4[\Qa3
M@KaXP8JTA^..9cBd=KTNa:De?d+?CdD)V3@g]+6HNcdXN7=5aD10g#/A(SgWJJ+
P7@ea4a:D+6V)Q7@R<4Z,[gIbXS.^?HeE-H>(N?Xf6P@M:eMG?5:;f>IXIPR:78e
g[a#775NQH3W(L(>H_2:U,\-:9b+#D+Qc6[YDAJ\7e,R;AWS;<=5J88J5:/YIf0L
H8AG1.H(B+&:(R.cXG6/-UbY+47bGLV>d\bM.EJG_9@^g77a\W.-6dc3D>DK,)5[
,_PGI[BIYP]_EVMZQC#OF=&E;0bPJU.H^&+,O8GM;DLZ?(-RZdDY3_BN)4\M5_@3
P6f87KcP,)4@+b^6g(ScZJ9P?LH>V]Ka.9NbSG3&8E8(]Z2Z=L2II/D(LZXJ;IUc
eVJ-.,ZAK5edUI;.e)bAd.YC5+eU(3\#f]<HPbJC#Ua^NYL2d.YK3Wb_/Vd[?0;4
Q1:@C.^;FT721=7WQQ9/^?-H#>QR.TL9O5eZF4(B0DGb[(>[:OWQIJ(T^J4JW[6H
S@\3NP)WNgUEf:.R\3b.Td\RI3U)R5gB@;>fL8N&Ta6\HREP];)(add-0]_X<6U:
e-(60)eFZ_gG#\N_Q39gC4eZBY#C)XJfSK\9<50=AQQCC@ZfP]W9B^:@ZKY1BYG/
WQb?Vd:ODIPC,&W8IYZeJPd^D54ZcLMfQ./2b0V]VCN>c)HRe2bRU#Gd3TQ:NK)M
04/Y2NfE2R0<fYSB.EcSB^cKN3HT;ADN_B5a=7KRUN?0SDaggTaT,Yf]b)6U=8/9
Tc8+B/H<=>fRR6JF57J##.\OK=S5@670e_R/LG8(Ea1Q=bZUQBPYT_.DD7T8;P5I
=6VM(DfKe,HX4W)@H9?;1Hc(K/fCDM:.D-GCR?Z=K-P>Hdd7;K/&1V;.&HI0O7D1
D>e)A:ZVW,/5fg?IQ;#]4#fNO1ULNE=ITCf+UC;b6/L-_IH[UTGE=MC9HJ:_<CLJ
L7F5855<3,WgF#dVMWM))X#8aE6IBI;W<I9O5SO\;A5=FI@:L)#AO[-?NBUf4U26
bMD9<LZFV=IL5(EZfWP&.2=g6_ge6AP4G18(F?B=+1e)/P>GFDNf(R(fTN(PSF0D
N5\DD37D(W[Q=a^c,-PAMf2LXKK0E6PEF5b;#2TAFDUSJYX,7-g^DAEG9,Z1K?gY
I(C+DX,g(OM9?U9R=O;H25#DHcZ0T1(f_Y_dTTW2@0FNU=35de\)eT#H9I&E:82A
BWF3ZRF?YCLJ<V2-Z_(Z5WMK?4?3?O3c59Q@:=<7>Z.JVJMUOOf8TAa^A6NfDWHO
]gEDb:7.DO4Y0[]=55/PW9+1M+5eRd37CRO@61BZf.S7[Rb#(/2#^_a4]=2XJLN<
P_V)Q_7g7_Q8=03-MgJ^,Y1,0a(DM<+U#cA\a5AWc+dFH0O>IO:_0)=c?3S(@DD?
L9&U.P8F_Q)6b@9]Z^0d;:Yb85RfK&M?FXB6Fe729-bgMED8:3-bEP0/Z\ObI+(L
d8R,0VV,B&3aeM2(Yc^g9_11Q#c?+28_,?Dd>a9K^,[\.Pd8(f<,=+aDC7IG8+&R
6Deg4?U3(X[A@5WOUPP>=(OZRU>dBTK;YPgZ&N6LW.T0S_,_9O-IO]BADD8T)WTM
H?C.G^K+PO=G9D?V:.>7/9ffLYFZ;+@g(9B-645MMTcBPV6#c3QYA/&1?b-GB6/9
1)W.\d8aafI6g(#<QB1FCI?f-bdAI4,.@ALD9Q-H+L@egWbF9VO0^g-6D:f?:;:+
L&1)c,-(^Hc)E_aXb+ceQ(@1U7IQXW9J,fQ;9fIHId_Q+>]+^M<a-e_gXSE2RN;D
?VLO&gS>>F;eW:[;K&Lc11?C;2C#+YQB:+7gP<L)C8.[NFJZ;UZaRNK\_eK0Lg>.
T9TM(3H#V7Q+.?[c:^a2QbJV&^fJL^CO3eJ&a-W]@C:FO]40TK,:g2@@(bG[T^0G
<[XREG[>F^Y<@d_C/6Ha(Vc-^d+e21_#[e;Sg4[?-(^=78><<YFI2^81S(L?)d,V
P+1)gO[F1&38PbLN]#^_QMMTc,eaG:DA2E,TG2V8.TJg9)LY+eg,NP;GH?^^.ATQ
4dc00/@CBL+^Y3+.BeRODS5#8QH9##<ASY9b-_G,AcF4);46;(;;>f[8W:12V5,M
A8@:9#J59-Z7QbZ\:#Y2WZE6QLSJ9>KC;/UIN&J@.dcCNI;<&/Y;9-@J9^..+bf1
-g/-6=&+(.9Y4NGHX[W-S\B)M&X)Y0XD3)f68YGa4b5S1[:X+F)eJ7,SOG:,c\B/
Wc5AP=)d@)X\-7b;2:a9,[;[=+B+)@,I95IM9^-G6Y,\.IID1PEHED7;9>R:<-NM
2?bR0_#BH((>\Af+fL#GY,5b8&USf_g21P5dabRLc\+\ZQ6=5FA@B_c:V(Q<@&?7
e>D<MRD,=d)/WU[,b-[a629TE8Y>O#OA-X:[?Y)UXP.5)KZS89?(X5T3.CaDd([C
APH4NVL]/g(WFde0dO4A>GDR3<7;bL/2b4,T:]^HDVFJOO36?()EbU.G<I)B5VX?
_59C01O+)L?>L.2\3YWf+B+D^/?b>8-E#BEbB;]5D4N@CUL^/J[aH7SJH4@<O2-N
aPT_==g]Q&_-P(?3A[OR]D()OL&,f/]E7:\,@]37J4P9de0#S9ASGXGMcg@d(dbT
(<2cHEH,&^[LA).O,#K[,GE>J>IL]NE=M[AIB=H6D(:g9(g7>gAU]?TKD5A31=H:
N5[Rd^.O&Y2&cTL.dUgL?BG>.6U1a+)7g0PgD-P-#Af5a&GXKS1+#e8/Q&Qd,7O=
a,@#4O^X=UMacIa1)dMUQb.E72I,b414V[WSOF(P14]CfdO5g?70_\RSM<c<Z@3W
g1Y5N>21V0@,cB8f\/?6e;?+M-Cg(ODQ(XP;]_\>)X9U7]&^TO[CC>.cgCRNeNb/
O4cHG##5IJ7LLGAQbIKI_KFPK3M0egQ[=,FgbPa9dS1[6>O-0/-ZF+HJWd_RA0:;
KXF15^[V46R5bY7E#e5WA+2WAg?Y;I(?99ZAT:LYEaL:2NSCc;B(3bKDG^A)&BM3
SG?2[Y)JT^c5*$
`endprotected
endmodule
