module DateMatrix (
  output [11:0] month,
  output [30:0] day
);

reg [11:0] month = {12'b0001, 12'b0010, 12'b0011, 12'b0100, 12'b0101, 12'b0110, 12'b0111, 12'b1000, 12'b1001, 12'b1010, 12'b1011, 12'b1100, };
reg [30:0] day = {31'b1111111111111111111111111111111, 31'b1111111111111111111111111111000, 31'b1111111111111111111111111111111, 31'b1111111111111111111111111111110, 31'b1111111111111111111111111111111, 31'b1111111111111111111111111111110, 31'b1111111111111111111111111111111, 31'b1111111111111111111111111111111, 31'b1111111111111111111111111111110, 31'b1111111111111111111111111111111, 31'b1111111111111111111111111111110, 31'b1111111111111111111111111111111, };

endmodule
