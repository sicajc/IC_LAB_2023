//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
dS5qaGwutD400syVOdUXRF8a403PrXLHN1f3J1kdD2W/Fob+CM/9nxtVRD997QOC
5+65g5Tkw55YQLSK5SmO2HZ+SKyjSeTNRGSQ9/CQFmN8S3xwjKs/wBqi4fwdY4y7
cWpFIY9zA2ARW4DToatDVd3Fndsc+tJsUDI3zRuYL1rlklCZUz5HmohMagCl4VAL
iOuQowQ8VVtYkCyBjUjHY3LvAnq63LU2mz3aTX1OxT4lnqhGaqJXTV1POCH2Fx8q
HMWJDGeWaJwzAO6izi+risLl8dSry91NN307+MVsGk/2b3W704JS/VMRoKDd5sbs
xWAV/slR3D3svi0c3YuMGA==
//pragma protect end_key_block
//pragma protect digest_block
1NChEH09bYrHaSTC6KjWZHl7Tis=
//pragma protect end_digest_block
//pragma protect data_block
KE3MS4JCbY1vFbvBUEjhoOzgr+NLPfbU0qyY1q/HzlmQa1CVUqPxaz5k00Gye+go
OFCeVptIEH6WXTVyFPaXubcFCApbbQIzzIaRlPFLPnajztXUAy4D1QLoWbpfLHO6
IfiZ+STJ06pKAEv2LHQna9DairGSBuiXRLDYSV0WtaA+CpLZcH8Fr0+r6ZOf5jWc
7b4mk1BKsRTKxDVqBPhqYZbpJAP2FRRCpA3kwzeh9LEPZlt0k8OXZDlGyLRTzeLb
vbevl1w7Ka18BWYdZBx4yaj+n+/PDeonoQWD4JmcUpXmBHIhCxSxUHnKsQUPaQSC
nva4EcOT4h1JVrcw6tr39Q==
//pragma protect end_data_block
//pragma protect digest_block
GFqtM7iwI7AlRJ+EAXS1jL6dphg=
//pragma protect end_digest_block
//pragma protect end_protected
`include "Usertype_BEV.sv"
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
pzLVBCHCw6FOcdXY0Xt5ZtTC9jOeFU5LQ3Mt6vbcH5GyAm4ejm+8I3nsZaTFEGI3
fqsHzAHcNln9bL2kK5TZNrVWlrM+F0q0J1121/lbvUKEaM7o4gaNxmEtsOoQRHZB
b/b93P1C8f+kIArGZpxHRhgPUn7N6tgetmpuzBiV6q4FQAOcuhC/H6U7GPI4TSaS
ZR9nEk/CFTpTTsBJpl3kcXE5cOiSJAVvkleQflHj8vXGibI6UoOj0JveLecu6sZH
YrxrpP9QrUnupiIOQNo/qVTit3wS+txWEcbn/l/pRDVv5lj2N7glSpT7WLuomP5p
pQ5mMcyGYjyLNRgLo/ClzQ==
//pragma protect end_key_block
//pragma protect digest_block
C8mrE5Iu/Nw9Yi7UKJEr0Oan/d0=
//pragma protect end_digest_block
//pragma protect data_block
2FJ0EmR/22hbuVYLMLPTUOWuIoYlocO9bDkaK5WLwFoxtYZXiGGeH6hTOJljEkpi
9SCWuoeyK26hJ07epHUj3QiGUf33bRe70hdaMRwFZqaFxuD2GMIcyL3DMRUDyuCb
Uf5yTi4FefSJKUECPnNFxs3vk2fldzs072TORcKCEbhgCz4ZWGGpw4UyccE4bPmU
kT34rOQIoKvjsBlNzO1FVXXOHMET/ihMR/NFCyQ+V4Vz4ToUvj7A4+FmoB4gSGck
Tp+wcXkrJuAQPNQSliePxsU8kZd2sbtNLUocMaGNnYXvC1AN8weUJR7zbGUxK+qG
KgGheZMUYabkHSrKy06ySqOULOC8xRFzYVPKsi8FWPfe5++Tkhq6C5isIxjamYEk
If/nMezMBuOLoo4aWIpURTMM2IAbxg2IVxZDfBaiVt9q94N8lmYpoPBSml3lNguw
l1/aLkxHV2Cay2im2KJlMwYr2IO+unczPPnxUuoQEfvaSWz9NrRM3k3JluXS9Hlj
yVOXkcLKeJnPPUGj/4HfeON5SuqhG026Jfk012T9OssopdZYEs1VyL9swQ+z9hkD
3+ztHKO/LpO8UlrpkgNEEM6LymFn8+2jscAOj+0d9jmSTA/yZ3S8nx6xa6xBnX6Y
QaFyE7Y7p6yuorLQhfpUQ639KspUdRXbUCWs7sRvGZrak55tMT5gaa8YRfN/Uc4m
XX+xDV+96kDETe68i6gw37ifyryuJNxJuhJhcz5CJW8R92JInyU793h990swg+tT
DqKqRa/y9o+0xTIdYQtiFfjXpak92qvqDBo8WzEMOXUw+TdhzGVQ+jqHNtl0BJg/
y15erSv1LC6PogytNApi865opNiz0MNGdGb72DPDmNasFtsWB5kRQTZ5DdigmAxo
5Mdf8zqw+MGV+VgLjvXoOzvlXttq5yKAH+ozZRa8xdYSK0ZJtVb/A5Pkgooacqoj
NQdjce5/AMin3bnVCB6vQ50tlYg0luIiG+1tvKxpYoCK7XlH498ne85aU6b3QGHc
ixHPdGZNP5HT8345zQ/+SD/PhGnwh/4fNQUhi2XipYZbRBtbQ7htOVL+G+Hg3fNO
y/oXCPiDc7WTlRLoqhHKv8eOs/QNzSCgSfw/1YUr4fdZ24LrnRnpMoBzcioj8t7U
wOTpaB5ppBHCNZ3UeMzso4yX1siFeD9LxelxkYYlIbx4TKjXALC0460qUa2a7NaL
7aTef9FYF+rZbp07uJ//QmEVgWBlfrQWbtUd0dJbGaArR23yFVJFWuHOo4maVuZG
RxCvUGUFtsMgBrWD0w7UvZLWntn9EUWanGFdxkFDWrXp9L8Y1IAlHonn35WvPLiG
DAuTDr/9PiK01892IWfkJyTO/wYNA4GtGndV3xlxOUWi2xdUDTVLrzOnGN0pvqTm
VQOg29+b69e/igGJq4b0jPGmXdds+VDK2O8tBZYDOo1F+I0Dv7UfypwnfUzQoETV
kq1qyDSh2g2UCWvRiFTKpyAMV2fmMBKxicoFyv4JygJiwTLVYWzNT7ip8sn7bNVy
qLjUjPyiCDZZyQv+vE2FC9m99K48cAXnhRnZz7+uYXTyEa8tGmedlPA4ZmUmNWwC
NqNokrnHQUToB7nyJu6JAoy51UQWuFRG48Uc09DU06LmJnusiHlET8TEFXN9vX1u
piiZOCd89F2VNerwg81gtqqm1ctkpD6imBIeKKIC24PcxFtsAg4lVX5KJcyJYovM
HFILqabQy9X5Avzuxf+erqh63QyyJcgoAJGuAbx7WQIob9k4beQ1SnWpkBM40HpS
0yOV8bkOmLJfZ9Mo1LmvsaFkD0wmiaJ70fO7TCCEUidyRJPso26Il/H0wEkBZHX6
iLOEs40rcFpzlkcSmhHrucV/ij0vUOYhQmWzhThigtfTGV3wonTbtkP7dDS6HrES
Uzn9Rp+5ogll571soGq04+3TwIRSY4vuJlH/neY0N8cVSKiDXhJEikCuBrUpn47/
rE8ZCrlHJWT4RzpmPdbvH0XLa023GeVp1ipEUWdC6mPPzZFcyzMid9zp7sHdhDwx
QQCvVANid+Ds2GXLXxpvaReJeGECa3CTenApUli9zfPlDdzQ45JCqqUSFCXjA2yq
0W4rYQVw+T6tJh44gL7CHawg5v7BcUVQ2Q54yHVtV81sB1SrDqKjbmj220Kb1b1N
O/GUGi1ChuaU6iniW2S4sATzNCEt0jZL/2YdzrQugImNTM5xwomYO1zpisdxSMXD
W1AJWqL9RzNo53hvBLqbZFmb/T4Muxtfd+odh0+kf3HPeHugwCU/It6W2oy9sYGN
jNwrttYbGTdkk7Psh74CescBn7S7BUU3YVkgYNVKuKOTlc7oclIjJ4ngHAf7xqSV
hUXP+E2C7L7ivWog9R7IJBOJOc/6sRri/sHqHPcVSt0hefhyj+hcvOCksEUdPE8I
zeJQBuHNBmL3v7/6xm+CfWBsotASRHnQgwDUR5/2JQ9ZNOgfl28cV7XhKslcBPrA
W2WUzYF064LaxNGzld3eS3WjVOnAt/tXTdedLgRTTj0Y+dneBVaHvU++xrCKmZer
Ux5r0gV+dnS4zx6xiZl5vjbFMWCgGcjJ4MwbzTHruGy57mpLY7rphpsHir/zuhK4
T+SAgiUg05zRH+QIuOBldD+sgZvQdQzMVIgrPznw+zaOV1Zu4BNdf06qJM8GiK7Q
caeeLA1DC89UW+fbGAUUVLbuJTH4eabZa6/k5m+Ldrl+HKppyEp8BfcqUZ9hpkO0
tL01XeHxJJHJ6XRQMWFhS2YL/sjEY1duICL6n1v2YsEoZWRn5AyOCXJ8KjggotQ4
ze+H0zVYLi33Td3aM9EZklfUvY1bMQ635dL7dZYuRlzO7FA5piw7HCPIJdKJjVdU
UnAfvgD6RhZ5q0ni3Kg6DVRy/gmvTT4Te6DTnG7Swu/C1VloTHMJosdoUqisUAwo
dOqNu0S0diAuCLmzUYc7z8UA/YTV0cBOGXRPlEFD9Xi2u+i04p7TPAHpGdvD4SQu
3FoJBkD5pbwBWzie90RLY6t3kQRiPNXWRY1L0vqjr1wVdrCQvtB2FdGxzBO7iZ3Z
3SUFML7uDbOt/ib0yOBRFcrUGQfLaaBJ83TEzAB22m4BOFihuaEHYKARPLxcav26
l6FSI/NWxCtIuPC7zE+aeWm2jh20gc6V2ObdXUkoye0XpT3Z7BgXuPc5WPqaDtvf
TLiHmwMyvQjJGHN2BQtTRQDW5BL5h9WfJlVJIaW00mMgPEJ3S0b2fsuZDAaxjqmD
hIFFc2h/IqYHKuRtsuVcBSBETz8eeObUw3BkiUMmAxdityQbUMh5zieGfbSEEmp2
2tooaTA3giGIUEtvk02/hcgrWB37FHADpqxVSAENsNRVPH5rL3DTiq9GG8RzldzR
8pYKygFpC5eILIEn6nnvJygoyqc4aO/I466It3jsxEwzMnG6jOkCudZsi8QPFmN5
aLKDOqXwQ4SkpcadjOcYbZaVmuFqOJ1Ghq9HKapAiOEddYaj3q9EUrJ/p6hWHWLk
h6I1fc19/CDL8ccW+6pSWS5OXiYx3CIVMED07liPsIfRtj/q7mjKSYd9iWLAKK2e
Itwyo9Fg8WTKiMFRe30rtrEW+SPklqFdbqLspLxEv4ENhHWRkdk52k+rBTtqoqmG
lle9qOyd3gzPDH6iyIiJxFPQIlpeWti1roc8yHox7+6+9CIEWRTg9bl6OgcuGppM
NhUatm7zLwM3lSlpzvB99Bmt+sjizLng+E6gevTW3Y1V1QhKWZm4EZ7ZHFnQOl9v
9W/OMDp7MjZ1xbHGlBivK7LTwouzTu/F0dfppsi4+E0XwXI/0R4nWrt9M8gThVhS
sAj7RUCRK3aeSmHxVIphsvdVKM+sitvLasCqhVHF4VGXO95vD4BSp2wXqh83O2jq
shwogHenK2Osiq0xk2U8OmdP9xvw7Y+kDGbJSMukSM19Lm6oxlEkdaMLz1tFVreg
Fd9zbZy6n3fBMjK/CKJ9UFlP42WIraE4mNWxBlut8j3VZ84hNCtostgg8wmYFe1x
L0QxeBbYvMoAMV3jWomk1qrXqgDNEiHtvrzx95nnXps18lW+Yfsqtw5lORz9LJnm
t+ARqUPaoy0IidMAeNuLKUZUgLRKhBO8JZpuR7H/ZJ0GEfgyuTjNcSLShJsAm7S8
7OvB6CQMTzZjDKzh+KAChkQotPZG13llLtjVlC74gdUyhTincT01nTG8xNkLSlJ8
qYU2AS6Y31Dw37STWlWdEdUqk1aGE6HARWHryEpqKmoAE2OebfKCKVpCd5GN4kl0
CEroOvTLAF0yRJhTkqi3E0lKE7Ajf1iu6PMTgQ4oWXeCilxIt5gUID6vRgmMTSV9
d4qqDkjAKYS7GrAEE1GPVuHEuT6yHwo5Ase9cU7zhmBjfkvqjcUUvXVNVsYDP+1g
CyZEhTjvtomfY4+NHZeqGW1f0goByZ+5YxyO5RwdhoaYIsMqELsskDtqMc//A3+O
/5vl8OSr3nNv63gkDuhv1CRmY+uYzoQXxHWfHHOJ2FoVrqYSyIkRcdA4h6Kh3L0C
TXcUsO2N4NfkdCLG6ISHEGyUgvhTHd+tbqCQqzGVMxP1klZdiC2s6MJYKN/6R5gt
4uYjevYmQmdir8/93FqL6XBU48ApJGYxTm04QiYafekjkZzXGa9fzaiM0ytRqLan
dp4bMqpSNMvGma/QPLsfpBXR0f2kyINabgtrAbGeHFOAH3ILTVucjHU/0uDESH0l
Is7wHfpCx/1NtOulHlQxrlALn2pNot5ZQy4UzhhtP4d3RAotOSAHtKxZkLbPGgLi
Z6bYXgQjwrUeoITfnCqE7DYQ02vng4Y8tQ4WqZwC/jhz1I1PKXPIIaVuOtoKr5NT
m3oJOky94OEjxzfQnuQlJptxjMR7Okb8zttsrfJk3JS1Cm5UKkzxSxU7Jl3VjZ+c
yj8MT8AzmqCWJVkdy/zcwl67m3DuG0uuG9CGoyG+b6N3m1j4zU8OsZNCVhyOX3E9
9Oa5JZmpMI112bDRMR2D1R6sCRZFy8R6/jeIvO5ku5hSdtmhtugapB+yvDgmJ+cN
425ZSvA4ELzQxObcBFFAVt+JYRhrg4SMx48OCGDfOaT96XmU26hpGWInNqfvt5fs
vIVj2XYXa577Aq84/ik7+JIZAsvQhuxRQv5BP/LQ8CgnOcPvkD60fyAmZnNGoTjf
nEMMKQz3oNwEtYvVKaSP/Ofi3N/SVLr5dccpBt8tP+hIEE6owsnxLzn43XXvffQB
bG2KGmKqetfhoJ8+Tv0rzYgCBncColFjplCI1tb+L03lO/mQXEEQ3ttQbF3/SSPa
zMqd/SBKSuSZUCDPtGNC/jZBe+g9JzZVdHwVSmpXDSBJTVAsuaGFX3UBTKf9m4tA
ApyWf3iHgwmGb26t0jnXlNUT0Xj/2/pfjUFTjRkpY++nVgScS9AsUfSHoeNmuGDG
d8UjCQT0h6njyU+6xr2UtMXc0NgoVftUuziywV5hqduXRpFWKAdsXjUjhK+z5L4H
oiz6YYAKKYXdsScLOdif4Y/Q+VMW+uwWKOFdoqg/ERQ16JUhsWHzuACUEdgxbdLz
V9F0hbf4rJPp2OG+uZTzZkbU6JIkpYvAlSNWvyKwFzQWHI0UAuU4GA03d3qMADK3
Bp22wKI1lnvbUlAQrTB+uwErRfCXyEVFTzNceQ9ELG+wRKXN5ePa3k9qJghSpWW9
zuUZ1+IoxOLkKq8/6qyKNQmq+Iv9CK7aytecWpE9OcqHac9oUSqP3xZkFZXBgNaF
NySL3vWv1AjWKgf2KGzO6XCgR6ik2PkoAPEWPnBGedbBwxGFBeF0OWJIKmky3i00
NLQi26ADHaMcLwg6NSCqrfAfPnHEv46F0TH7OYrCNp3xcHXkvL1iaWhtpxqbWxZN
vK0R7c+UBybcbFNL+aZp37TOVRxRCG+PrlSnl/xIK/1tSbSoN4Fbkqwg3LjSnFFg
OYlTRIkrYe9qZ6QHKsFvFMvqycq4NzVy5Dk9pZsRXDC2TpeJ+Qg8yzW/GEcQbOL2
NT1EyuO2WnPL3Pbq9ndmvE/urO34KKlnzK9JCKYvMoHSFJXCn9jWhZVmsbaMu+cY
F3N+15v7JHDUtFSIVlCQ+6qdOSZpUCpHSSLrHAtfpWLNsAhEbkAzDJ7lbJLSdBQv
BpkD8xzyuodRsZ5NU59kKciZgu83ib9IIVe2/bFuo3lwvsTN0IL+qQmvF5GwyKnL
/fJ0mHOg86Sl4Fo9vJTMHPY7MafzxMb46nAazP4oj5egqDFaCdSLw4/YAztvJWPm
HopZQuAdfx0J0RbRAdWGrk0MlGvfJjJ8UtxcmKQUh+PaUnRyGTTK58HAo0w8C76l
G3v8k/LFzEFfIExM5A41ttMucODbOcsQcHt4+1zcvNOq8PuZK+1NgRHjfCNYC/Rn
R9QtHrCmCviEi+p0IuyiAaTP+2OVeg/AAm7LR12357qVwlTLzS5AaNyUH8Ms36EK
e7KQGFcMQ7/lKTqeaRqh87SioceBi2FikFYJ7y+aZ+uOB3uwyMvmtRmFEluq8EUd
uUO60B/4z3rSj9EcQion6lsqsrJYHJtCK0MQrGSf6eAZFnPe5TawZACs9bDMzJ/s
I3jaFATxEsNhCnB0jvbGeoU4844MYmLxEVR2PYRALJOiGhuvK5mNIfP7YLAaBORM
am0Zz/T7fwQ7eWk3PPbOL2yGYF+AsbbWYMJp3tIJkx+cCba4VxtY/KNuHmWq+Ymg
jDu5SQZO3yIA23kh3N835Az2ll0CG0za23fAcgNL9qiZtz6he2KcfBUz7Kwbn9j7
JaWZxmeKfaU7ALq5rjZdZv/C7SwwZE5N7fE4LnPOt77Q1XeuZzWRU4vH8/hqrFWm
mRLX8anLSXk9koYb7HQnSej6hVbpOBo6hP86rzkE5bZvBg2lq5fLtm3mqPPKXKko
lNP9lxHADhEtKeoMbGUR7jn6pWBdhdcD7HPCTKYIZd0GBMVVAurvvo+Fw06a0Whr
hu49FpC9GjtpibuMXgys5nOrnULkL66SjBaPQ/zTTWhUvmMKEI8Qg1MrCLcgz4Tt
j0UrHvRvIvOH72GeHXDID1T5UgN/L2uAlQ8XxmHf6AUqIuOnToWqFJI5gH3pqJRX
1FZXChLnDwww9/SxarOe5k8cH5pkWC3EQxjtROKSb/4r0QY2FX6OrSZP0F3sytLV
ETM+AV5Ht0/+lhaZ9WbhqIFY95uMdpwXclmWrkakJexN5RCWrI09F5d6/tsLM+lw
ndyQpKXD4cm3ofdCpwE9SZo7fHA/Da7na/0ufDaCuHFqNXn5eSYa8IVgDIbGrVcW
pz+GECOWXcG+cSeOFuHOtioayRkgwUNrctpR+tU1B0Zg6fcxRzc7+hUWbQqWpC7/
FLjgZpf+7EcxNndY/S1J1dgc3eWLkq65ghdzQ9seH1xyEWK0nokfDE/eHLwOvwcB
YjD1P4GbQ/Wqslp8NJ+LzLZ7nS3SX6WnlmE8te3vIGbXfLaM+3zmzsecbSIbszAi
EYafVqLzJwBlWDrF4jFzC9QOhdbjQkEDB/7p8DtN1EXaGCAMgYKlgwzai/ufeAOm
8FcXMZ9aAgibgmwwQFSKIxBxTgxvCDZJoJTkgXYTpnl6tABcnNl9Od367LH1Dsqh
lbHaerLDBIaf053RXDKpCMx+rJ+fiCVzNWUCdJOYxUVFx8dkTABZ/9AV3S2c6N35
r4SEaDJk4N5uhUlMVVpLOFFmB9dtsjJBTOPWiKH1eRrVHpEBdzIS5hzZzi2rAwBq
WsuWIpSG7pKz2qvNaV7E+5xlaLHSs1dg9u3l+34GHGSpeDE0pnDN3iVWF5uwPfnM
7nmsokxzAiOloDZovM5L9i8dlfCZEFKdyVwT2Qe7cxZQFdyksONwy1FWsg1zKswE
iBLrrvz8A/Jy25uMJ4dtVPAFMEFq3+h1GLZCcOXcdt4cipr3vF1mqm81U5b2OlT9
hgVVN2rEx7/SrrI6tTbo/dLcWuvp4SmowOscHhHm6ivb7NV+BFbW/FcRCeAbF5Cj
HHvF0Y5/5rmz1igbFVIyCo3gFvZ1k5rEK7Gsc9p5R4CnqlAtIcHt83MIf9HrEH8n
kttvdd/fX0Zz1POMLF5YxbCnG1NCQcz/+34qho+WLs9Z0zhqKfVswzQD11al97oe
7EEK87r8fVcbmeyinxzEi/ND6Jgv7CZT6nyQT820nT0mr0XAwrMlLPpB4dNJ+JKD
mtThE2R7+G9DmmZmmwwmdlKvBW6IlciTDgAOIiUOOzxAGYG/0EjJY9Mrq2GCE1VP
H8vWp58quMuVIRaJ8lST1/5BrMhXYK/IfB+e/s1fYlQ2VbkzG3OEIf0zOb8DpSad
HC01TBhSBAAezdoMuyhUtlolzALjeFthT28VSU3+ybV5V8PQIBliqsA+ahn4Luhv
vAmXizPFcDZvUtlOMmypljJ5hb8aIs/0PTzIQqF4idKPqatOAGNTXj61m/7t+lFf
P+lJqT8mcdcDnlKpkbDUlN/Ks5LKmZxQmz+ePDWim63olU4UTsD+H17z3L4CeCOe
nbbQfNkwOC0Hm4kDRgHNi6JN8s1+RkkFAvKZeUBet0EpchQz7SfoUCKpjzhxf2y9
5+xx6ruPKAHtHQ7Cqkxmuxh/+GNvx7dUCn3l/tOAToJg3/FUyKOSshCptOpJ15oJ
NAqvKkFdFLFlVtquvoitzCh14skFgmlwN9/psr+OuCY5BKhdoZaPnejyrGQCEWtj
dDu3Y0xi6G/RARqCO8fk32PEZl/JKMnbM8rhJ3eyp6ToIK3XArVyZ2ojmAqSH+oc
nPz+2f9lA+31hJp9Fh3vUmq5264/lSESgyZ/+oKaAkiCK6TQkaD6zCaC2xVAUxc5
zARmIvmYhk968dEoApj+LiRmRXXbop1Qlbf0+cCeaP8Zpr3hnPAqNkFEAOx7nzL3
c8tGs+idb9I30wzWjfe4W9cUEe6qE+VrPJuuHb8HrwDudolSKgvmKE+P4FPte9jY
3AFGuft/ZyIWOCNxHgh9zFGWwoKfMydHQDWh1SFVUwsgd4eQAswmHBd1P2zRrK/Y
g/rDYzwPdpL9+ejaRjX4CE4otWjNGklNwaYPMcp5rDzwVl1remMmkbBHASqlQ51K
XtBM+xk/n7mZKLIUznpx/Oi7zBKqoCQK4+lwLRl8G/A9MRtgwviZbMjTMnHHjShd
xAcN3W5MUS4kQfPC9qFVptQ0C7bzJCDZoATXsDdD/MrfJ9J9JiDt/83OoB2jpozi
xjYmf7NYRvjBZdyQ1JlRo9ExTVw4ot95hRH+PkUmsTjSU0qoEPfXvaBqFeEYMhrr
RFVSaZx8KUmiSvxs+FUyjY7eU43Yl00xF2ZjZldK1TudXpkT49+eWomcDJgwGO3Y
bvv11FUA369FusFht4QTEC6nCboueZUvteN5J7ocA9JXdhBrqvJzk0bFs9K6J1JN
hksXXEFqVa9cUEmiZnWJVsmitgcfjqMFCVhSJZtcesLUXs5eh0S5BEj0CPh/3/YK
r8S1RHUMpxaOrlktWgjRaHd5vjF9Br2f+yY3Cxjl0Hq86QdZOTtLEj/8TwH0mR7Y
G5LfKI6RYrRIlVZJ7OBRa52FVWqEgGm1Uc1pDouiT/ZEUBjr9fXkb9981x2xw9Sm
OgwY12T0qKGvSaBInbDU17JtsKKUpv/ydS49S8uj8gBQB8a5cP/9HoKaV9E0r5nT
5j7JeKLZVbjjD6Gav/oMwNLlIrwv45Hn8iL3ps+NkDM4oRTVtKaOfMATJPrBFqyw
avtkxjSpIHNlV1G47CNEtxELy6S0qYznOOyvN16f1tElfH5EkvdgDy2Gajs1NWhY
vYcKGko/9OiqMgC5joQ6M89Y4uVI/ww0McreXerQV1QXazIcT+4ojRYTXQ7iXMJB
f4Nr1gsigAD9kaGAkkZG+4lyh2erxpZKiCzeXUGjSvpdPRmghhJIDmId5EA41bgY
rFLYUNv6MFqySM3SrFqKEL9FeXpFwIEWS2frsLo9bqXf1Cv2yVOoBlYSPNuJ7WWi
1ao9UHbRyabpKVUdhwg4HSEDaTWlxbvFiUfcybqOGMPZrqBLXnQtlC00NxqMzBWb
zMjDwtBYQqPK2o9OKDcyIXLyEoMICUxS28+uVCy6r4DgF6bIM8mPp/7PeuCmmk6X
Du4PE3CBjJ031tMGz2VkKObZz/168JkuEN7KnUjRmEuIYRsCYQKG0CxaCUqcSL8c
bcdnzFUVsNZivtzCLJr2Si1nfTvT7yNUeL9C5y5YsKjLToFdehB8N1c3U9WONjQZ
EO/OtWX5+EZwH6edJyNjcLSRRlqP7u2vCM/BYzJgvoZZODBN+SVIXrhKNLb3SiaM
aNeejf9JNOvnd3FZPE3/I9mrlcvTNKcfcwlHJIEVijZMycEvgl7OOaC5fy4WM0GE
Y1Q58TpzWElQPmmnu9LLwgYto3iKhslmRHcsVniqAb4gyq3Z5uE2upXllXyFPzSd
26I1FQXPJOkYYetYOl/VmbazQxd4DxxB4Ij00sb3nGYJemFrYo5OIV4HZTZpOCt+
EizJAm57C1JmlWewVqBd9TgtSWPZxtShRTYVfqDG0elCz5hy56JIZyIjF0p2gXoK
af+NorhNZyNg5YWR+VXAGU0t1zGqYIyFhWVUedO1WefQKzHVJlGLn1cjwPWB2DCt
kLq/9GOEEtJmAF2P1ggyuTSYMTL6kvsxqqbRwXX+p4kgfSPS2asmpM5So5FtUzcW
s9dWJb2maomukZAgO5v3NAnj9eE4U3ELsRZZ2+6S6CAsdM2J38a7dSzJ1A5ZFdp/
auOW+PbNN3zGhxzzm+JmMVl8LdgpNOHBxTIgHCP6BAh6iw8kYaCIJpCqDu+WWI9J
KZqq/ZSugqiRCINgB67X3Hz5GSLQB6TDiT8bQR6F4lEZ3RJYLP0R+tykqXGUJ/wJ
Of7xbEhDqghqAG2qDu/D+n7SnNKk0vYnqzuOX70J4BFjifyMrawjEDrxhk43U3sX
Rv6hQihJyvPxUUSv7x7QBl2FnWCNZFF9f3Vvl2ADhizgSsW3xqWZBSuUfTE4PCUC
Yib3OoCDDf9CRv95Zd2QomdAJyNLjVj0v35pC9vlAtplspBXQFqw2rzx0rOLrqpO
naHXEPuaZSX7rtTIgTki38C51fmPfaCQpJKxop0lw73yNsllsc1RMaPtkp/8ibxW
e80460NeCPGkQKyzh3mNhV9TePo50JpiID+8YulZGNnSLCHEofg07jCfaXUCeg+8
NQyV5RFFsCtiKxHwq25RieIZVNe7T1RZlH8ZogLnEMve3IEre0i8WE7I5/N9BhEL
kZTU4gx3gOr/Ul8lM+CxHCRRhMPNbymWAV/4qLmzzyLjWEcju18Rab7N2QPdX4pD
xzOGeBA5n3iKkBrfLakbd0hb4DXDgnQVa1avgKnRDy8BrxpRgp8kkvBloD1CD7BK
LmsXgJDXUgAK3Lbvp9cIiimhlvmGQ1aHq16XWoJECuDKLKPFS0wwfwkKk+YjDHdH
TdKZjxOnO23ShyuxhGXP7Lar5ofyjzFRU3VYhI9BDjl5XU9yrpxCyJfAJFLJvU5S
gsHmY/0RRU1huqym4R9GQmSvpPeJyWswvZECY4YqbYpk9lRTWPnVeLJ+l0hUgl04
vFbQoxtJk4AgccDKslg+amqBLjD7CLO5Dh/LEQ3679xQBYXZVnhMaOAwYHTWB0gi
4T16FwRYZolQPybmvZwRxFelzsnAVO7QtUIAgvo62LZz+r0Y/1ym89rMzHnnogJI
cLdIHm3Mo5c4uwhfoO5a5nckaEwJbXs7IHnnsIMHbrAspi6xePnIG9Ua5RT46ikg
sD1wOw4wAqvm6uif/h+mZ+al5BVydfbvrSh6ZusQZ08PNypL9wDmVYR64qHlOyaA
CHdO3+J+tyMfHhFg1nTjdVxydljiytW0rjeYRd51mJ2dcBwdjgptuB6T+EBTHHMZ
DWOwjk5Kk8MTsLInxXXEyTorlQ5VIQJCTfPOSdEzYjD+kqGpdW0MTNC7yA831TxX
r7svGE+bz2+psl3vuJ+7vuLeunR10lE9j+R8U/sH2cfknO6yj36wvjjzJUJgHYQS
q+mz+W/xwx6mGgalXatwblvSYVBxBgWAd2x0YbthWQmVTFtDgirV1T/ha/aNQvSv
l6dvRD20gYBAzEG01RB7EM76G5VPXrjEZD6cqeW/tvO50n1a+UkmWdGScnj65CDQ
cKMupZp1eTFXba7qvyOAiQLZR8a7QmoeInzGrymMsTlw75r6Pb3Qix6/4GXMSi5I
F8omhLKYHMrPkOqiu0c8BkmFk03PvTIx1BHWy1tWnHZEyLqQJXNJ4D7BXxeoD6NK
vX3U/f9kiKfmaUHhHMiSdmBQZn+yVpT8OpRsDLoM/970tERsOjhJKiC0Cb805NKN
jOhpwjOeA+9ijdQ935wxIR0TwrT/ghm/nHH+7fl8XasIyQfaNNQbD4Ug8BDxronH
iIlICI1KGeoAraUyzV51BvGOUEUqwpijhY0EjHYrGjKmiS6HBTHzE4wPhOGXTRlW
FVbnw0MGUwhWfwny6zhJykNDQmv0VKVgZvkLShgPdYhRwGWZC6/iz0NLhDF7SJNH
oEgrfW5Cr0eKH3GrgHzwMyLGfKgsDwoOz5cc3JS4dOxWUa95anJrDyjQOzGaDErV
onvE+0IKl0VNgXq/ber6scgEFSf6NAWA8yAprxudAJ8nBfxS9lIR31qq43AqX5WR
dHgo4P3QbeRQKnpD1+Fj3Mx/GJ9/eSLdqfDo4hMvlKotlrf374VXp+yR2NzriDnJ
6inEujbGeDf7bxbi/gwjEGqFvRqNM8YBWa4yfN4VORUhDI28Ypa+35VJmzjHbEjl
or3U/XypdoLa5KJpSRMkd3nPCyQNnaYD5Wp10IivXwrntH05rPkmxXvknXo3KpTD
OTep2XopetxW9QpnpVRy53NYsHePCVEYpmeNhKIV1XteWx7EyLOpv6wakSH6Vsk7
tjfL3s0CSCoRhL4FL+EPIEIr3tZ482m7Niwg5bnpwTGuyQ1g0fZ4kphhDHF3gJ1D
UZNmSdbR3m6w3KE8FO36UJruHQqdPvMQy9HTz9sTJZcfB5pGP562R+5L2hf8ajum
0C3J93E+0OaEOmkvwHj3M36TDESz/pE13cPv+0HfzOyyjnf1r0OC2dpFSnyJgroG
fxwFkUzBTQXG1SOWHaL5r4HslS9oQrMSItq3YmM0vdqkkY990vYPLu1+Z/CawhYt
+BTL4NxEUbYMzwyACMw9G6BVCVOLzdT7POt5QHmvZ1g1BzoI6vqdTHmd6oyffsEL
DI5mlr2qnpuDcSrmlGRKsH0qfJFZip80pCd0qAaF3mQdx/PVb7GldBA9AX44ZuSg
QCH7s19hypvZUW473byk4g4suuslt2qT9aMF0A5qb9OS2oK7OdgKNhmAAqvHICon
Gdut6i4WQyd1FL6DdFhVgtt5nWwfaePeZMMlUzG9DkS5R6VAAsCGuQe4V2lV+x9N
hNk+QUFan8xelFuOrmuEGcerS5DDT7Kv4zFZNrNMw82zqNN9Ra7xuMr0dU/lGYW0
yknArQhVcrKpMNhCP8SGoAXqwKUce8KByc2sapVDV+H3TZaVy+e3nKaaEIrvm/R8
2tfq1nonj2M8hYGzy1hUSeg++bFr7V+ziFn2yuZkPlRgq/0ZGhLt5cySlh38bZzW
sw+bByMxDRp3TE8ZNmLuuY5T9+T/okMcTgJYSBVp5RGZ91sVtfUmF2xqx9YPKbf4
etJ+hOhccIH/I+3Ia34f6q6BQJuENYV/M/qtKJ0p7bIYOuxCFu6uL9ufrSRPAPJf
ne6r6Xd7T2M1Xji5ha7nonPBNFivzVRHN5uEFUzOwSf0TTdBaz6enPi+QhSjI3ne
yJeSa1bOqnM0eiHl/j/1CdtjcecY5jjjvEy+1dlnrM76NYQn7df1rJGqSfYgTxMY
7/b2X80v06t5V9pvxFGvwsTG+7oWcqnYy2tHLVpqwiewFujK+4gdLE3gjEQ4uYWY
dDossO2ryR+VRz/3TTfFkfYA7k8WEfnokHuLG0Xji5zuFrX+LtEAprGr+fEfz1n5
8czKoecg/R0VY629gCgRjhjul/5ii8FwmTVuRENqK5dZzOjiKodDCsIqWZKx0vjJ
n6HiPEanILpmGlLxmPSGUhtSiHuzJDtFV7+IWll+xu8S0GznALSE15K9mX1BOfwR
DzpwQUnhasOg8Tq7RhAu6a3EwNIqF2q1X6kToe29pGZGQ4wYVr+GO8e2ci2bkJyj
9TtT5nUzhRIFaiYNWHNF3iMPMTPnfQsWnJI8Y0+fZapPYIazcrM92r3pn3A7UBEi
/V/H/wqpdApJ/YSNNw01GBT2GQdcGaAJS2n6NCrKALJP4yUfUifzgKBiZni3s173
NpC3t+dxq0GI+R+pe3FL30h/uQkOSgEiFWPDGSFMiP0YgwBLwCxm1m1wEwfmsrJj
vQYx18+CROjO5lVaY9z/JJD7IcS4k0eLXRKC2bLN09FrwUBkjvVS28EQsFP22pVV
LYwY8CY2kx2wUMBL2+RiLazvmm5w85gomrNALq+F1UQaSMpYU6QYYZ6ZW+hBdf1q
KNLoHtmVp+kFZXLy4LrcYnkL/z40WfpU0gBts9q3IeBbBigGu8lvh2nAmpT3qrFv
6YUGKGqwterQebcOsZHJQIqJcMMEzNB0VPo22vxDsI3VZf76pc1N4eHPRQ+Ti0DH
wUmtvJiQ2rCFaXhfvPk0PRg7Z+QF/BkAnMPkNZZhP/qsAvatNByvTwFOIf939orj
7ks3Ran9CpGZxXBDDr+HHE9AoBDAdO8ycfvpTrVCthvjBHIqLIj7TcnggTTS/CSb
LULzQ/kYDEHgIYPPL0+bBfXHwuA1JYc8pxhzLOh+T99H9bAfndNRCwDzdhNjvvDy
frH7k4K+i0g2wz+pDI6oF2P5rcxYLKbsP58PIK5Mhd8emGis43RI3Rwu6ySCyNEl
/bogf+fHQgNc4OCcjlIVQGRAgpQ4MX5XIONa6GpcBjo5HWsyWyBJAv32YQVburkH
2t3pzniWfVWN00JQ/SUCzCC41b8xJN1YCcL6echSjEv5EWYtFEEXbxGfl4VW9JGc
4c417lATS1z9PyL9xRagytoNn1H/+KBMC/W8ZCZQ2tQTjOsWEFTSXaoYpz8TlyQh
K1dStSo/NOE2oWg1GIQYnARBfiqx4lfpTG9ql9JJyQ+Z0N0yGN4QZp9yU+2rRP/G
RsEw7ukeDB+6Tvhjmdvr28DajOH51AYaoYpcbdOTE7eOU2J6DM520kpQalDMn/aY
m59qpJJVUaWm6ihJMYvUf/0BOpVAxmnXr2YtRxcT2miMv4o8tXzm+0we5CrCdQAY
DTQizIj1NMy4sUTKxLtwt2QQAu8WjS4ThSn+rQXO5DTQeqb/jycPIwBJ6vmu+ZLe
N4G3kpTN9lp1WYpEpRJ1R0pkJlO4CGZWwWgC3vaG1JhLL+/nim5Av4/pMdzDg/E5
R5dtDDJGQ7ZAfeSOVLMj+TkCfyDWAG+g3ajiidSyYm6t4k68apa/WLSreW5FoIoY
PAGnoisvp1TAJijcBsGKuKTryGqpTuigAT9q0WLc4OCYrOAaxpQdm4hVvlIfFjd4
p4Ia+UwH18mYsfuPvnTI9IW7S3mCrMRrVcRKbkdUMIlzB1nmvVXYiFL5zy5ACAHj
fhSbk+yf0ySC7aFaRyRbj6gXEVRrlb/NGjqFJ4P0KaqQB9mTmRF1F2w31+d7H7z7
iWOheuHmBUIl2LmKDsbvveJuw4pQeHcCqO8ATiP9eZrEXPB8xbMPqCsFZZMgW6zS
VwnGs1Xlj+unzsFHYkXhh4iaa123XT6bYbDoTEJ+CE4+7L2GRJkBYccjiEhplWP4
jj/Yo14zxUhYHVz/DCshhMsrw1HoI7YHXuFfnJDwp+RqHvuvA8t4pQJhGWt+c5LH
AEYNwuZ36/YRBeIbZxM8AzEiYrcVd/qUJwavAHhDc7KyLEbDKz7RMI9Kt5RGDUVd
DmxmxeMvUuK/7NbBzPaQt4EDJb94oQqOcYLymCzwFG1ucJNnX42i8VA0wLrEmKeI
fjbhU8SWIbw2OzwC8NvMOitHyrbC0NoKSu9vw+A/wAuS57IIGqjXQzh5sX9DAbT/
OWgi7ZI7rXtQGwTSh8s2JUeyzw9AjtUuQhLSgh6Gu5gYLcJTuhKe4JZHG8Aem31c
ODqK76EYka0lNINfYDAJuFQWMNx1SwuKJBifR9U5Fux2sJl+/8JxvdmsAwnpqyx6
d5ZAsUjpCiGm812ru0AdWU8Kkjj95AhTB9YtJaCxCyb8UzDkJQQ/Jj2cUELnHDEx
7zczVm1rDjuhdwWPSYXM9xDQV2z+Va3QBRJ8xA3RjsoiMAU3hCfK18KcAm3PdYfD
Hdd/iuTvL5VabTxQ0CGcmrB6i27hk8+yoGeVKOJJtjXynjvj3uK6Ui3Lb8tVgD16
NL8GoSCsaN73HZPUNeL8dqbmsQsowL4U5Cxs+HngaH7E6dH9NHEOlodT2tEoB/Fs
R/5YcYZ9XlnzNoDES6YFxgzdpF1pwtQDrtXHh63sC5cPL23jQR9Ncn9eQD4c4rMR
eh/CYOQYAHV8eCs37dMl6eJBo0kEhdUiNu1o+VZsh+ALFd0aCRlrVIzzZyzXE+fS
Nty6LilscOPZ9sJuVT6w9BT6lCukQfkc/6VdSkfdHz+ugNVhV32AATSaEulDnn1m
mzXJ/DICyrLcdzoyhDijOIBuK+H7f7ICA6iZivbkBHtffUJHGHNVBndGqb7d+Mg0
Lal6eikRlQXrRu4AwN8FjbLngYTh9Q1N7u5bYWswcU5+GDIpbGThRPcLZuKcDzCI
spToMLeTqmmvYefDBqw5h1CoQYSCf26FvZhKDOTWOgvINvK2V9bU7bmK9UzZt3Is
mfIJdpGjczXqAiVUEOS18VwPrtEtYuozJ6pTG+BDDMrmRl0h2fiZGcSui3KyR4pJ
ZBC3wjd2FrrQq8EyqGpWKQHj/+xuaIKTpwp3S2oZTdU5YG53VEvPImxnMKWIyCT4
c3L486V2dLGtJ+WT83TtD5DZjTA657/VWarjWt6hg5GBVagA0atjW/zvumVu1TIa
dSQK5lVJuflxLNVYY1CRo/VNAK55yKrVrZ+o7QczhvAo5AKKu4jUuYQgsouvWTdP
hAWkt6cFlXWd5jc9psxXh2CIazAgpT6+5yYiwNijcH6sbWXKoRIKwRAaQEcuD6OM
nMlcnKISATP2gKnIQe+K3z+g5lcx0eLAd0j8I6qqQFETUrAJYlas96buZ3KZT/GY
YiMUp4olzF8FrhxrMFmN+DtKVLSKzSGFteGbeHF3TU+qTD3qGRW1BDptyYyQyVnY
cd4zfFNjFmNe7URFoXk3VDg8LTzCFD+HyjrmenElPMxkXyHzZBJrBa2N2uUMr0O3
e4mQsXmYnos7cB3+jv4gZkcOcmhAWa5brw2Y+y+lMqmoEg/OLLVzMEAWNK081mUv
Xb2F5bSSfF0OCjfSXC3ICedngb9fpIPMDVFJtpD6phVUQZ6DDSs4fKvYYUwTc5sA
yRWpGyFsrEFR1ak+uU9UXZ0718D7NatdrHpcXnOEqpzx0POUaCzAWbpVkvdzaAny
UPnNdcA48Dz4P8GHEw4vETvmZwy7wKCeL8rACGDoNrJ5rik+KoWvN53GPoYdvF4Q
8VrSPa589ABjMh3GtvdJ3OEhukXC1dUZ4wc2geeZO0M47gtnwt7S49I2rvpjw9io
4R3huqgB14f/ah0uZr6EZG4XKNKVwJ918J3usNWEt5TUaTyuPAIQciraOcuxi9XN
zG2SF7XM6JmNyEFPRIzj/HlJU4/3JPn99pzZQYs82LU2LcaGn9N2bf0Gnk0xOWWY
QHkHOx7TjRcBboD2+MEv7/jFVI0a0yCfHRDAlcuOzMw5uzs17E34u5bW8bhhqbg6
ubqa8sGlzlcLKyRUln7WtsqZHliO9FMVKk3qamK3FpvfAn044JIbuFCt3ixdLIkP
afE9DulsdV+vR7tc9O0Ia8zb/5vTCkc043UbgQSEMgxIWIuJ+agFxAr5JvPYMs5+
BC/l/KCncgWtYJrdXEsdfZ9Xq3IRW+XPEf/QjOG5d8jPc0OMKK1NgcSv7z+zNcbL
e3guK/Qx4AYcsFEPO6iN6q8L3XW+jtY9tmfcy1AHNEQc5W2y4/0+pKQzKAz3pavB
WBtEIIWPwwcKFYqhl53OWpTfihFhIU/pzjVC8+q+gDgDPh38/NHLEgjl02AvCMAL
sNtu/7jwoB54brGE6wLMjVCCQdNpv8tumiyLxrewNwTeMGPkA62AzbfLBPz56mHv
9bDHyE/jy2MHViEmx1yZa5nhEfK9XDqlw0CqpvjhMlv3dx6IQ7Pt/HSvwsThB9Vq
Gw91YFd16ZOH5E5m4p8JNoIB7qdOpixCggtWUur3GoEYb4mvZwAVELFBVukG7qTe
VdwCZQblFbP11oZPZRhcJUrqm8as1302ddpvUhovNJF/rrVxy1NsiqweXmnxYyJ6
8IJMNGQWZktm4wjvdd80O4cdMhJ6LBa36JkYH/y8HcdSeJptFfqE+2X3R2CsCUNG
f3MgMhQ4Ww25jF3s++E0VrX//ipW9cZMv+4bg8vLzz4NUGW/6lxAbvgMGfbGAj/e
cp8GP+mBWQduGliOsKw8+vIiTz3OYOtpFap16FLw9s+ZEkYnik/XlOoyWldyKd8h
WLFWwDTDVqB/cHg5HxOgjH2QxUghX2MvLVZyZUBnhF4bVOc4UiGml+2E+521fYKw
wCfASpA1R3dNto7p3Y/f4ptTbCRfcM4MTRXfEWzPcdWHjXPfJB+FLQ1lCYvsV/ah
fQxy2BSD7yaJ6CqqZZ4Dcc87/S3eHSw27p2wcX/H2avDSbsS1xFFcSbNlkVIlf5P
jWKPwSjIAr7h4qvbYYd/j4+q3qm7aGCAaajw75oCriE0fKOvHK1DM0lsSGrwG20n
vSUImfj7q8BvDjfwzHqPJcjV0uKZS0R9vejkwYqnbAZgX/OSf/V49N7Ggjy5/fTX
jzBsKBVe2Bjdd+Q3cu/utyBtVM+TEmQNT+BtpiWaBDWsB+21JzZFCyHfaPqNqoJq
9XYSPKYwBYvhI/E518e/vQR129boqpHSWNloQENd5NKYppO1atHxwqfgkg4La8pP
HlTe1hhpop//pHYin1/iRPQRkZ1oEYabbWIYyPJ9tx6Cql8qjsfKhcALfGn6IPIx
vzgJRWkqaC+umNX6ZjbKszc9vmVneDbuyEB5SlM+++Ynlpgm0TrvTpybIEOqZO8k
8pQ70oEY4qurnhYAU2dDIdPYz1IkQwxiWyhpIWNcARGv381cwl3y5Sle4oWXZO6a
G23lkNd0pMD++/tPOFJXSjX/PMWwcAjJ/bgmH7pBRp19O254MMbVbMuROFAJXYZx
cbiqCQw5p0qQmgqKrF74z0IEUueRcJOqhCajwjr5REGa6IzJsdEhr/rvCJFai5AW
iajnKGOyQOZW2q3XwdXwmxLpz/TB0x7OoVtSvqcZYxRBJKgsqWJgNfEP9pWA6/Mz
RelZbTbhlCWPYsk7lMgcYuYZy2/Z/iiCNRyWgdZTDfZ2ESxFDqwYIW0GUm9TVzQM
RN0metYLefGzDK21bmVnmM9vrp2c1edtBESp1CDdI86UWJdQGr+SqZd12tqrgPxS
C5gaiOJ3yvfSFa4WLCxdze7oSUkbCQ9irM+8AwA3aFt/I2gA68dQ2FoUc0ibfkEj
ggQtmchjvXjIfVIUD6+ncAGvcVXHm0kB0QQbIV8s196PMH4CfYe5i8vPKUjZ7W65
myCEhNjl97oOg5EeejAv0t86bWtGAn3d2N+VJxCz/UHe900ktYtwbyn7gyqxJsw6
H0xUg+bx7FIgae9kzpo+iMHr1q0sL/+f0eLhcFL4HrRSHUrB0dQiNx3Edw4JRlnT
AHOm0THTSZRxaxphHVVLfanFzubtwBaBIo1aN1m+E9HaUZ0vpq+WgP/TAhzpJHxF
Y8Wa76UiaU+ZkHn8KlXmA7GnOr8/GZlqtVOta2po9rpIVK29EWe6wpENhtHUOgmD
LzlUpyP8pPFcBgLiaMyr9jT6yWiVzGClzSMD2IvkTJFxKZnJjyyA3E48jgyb0ETG
M280ILzfTTzqoEYugpo5h05ew562C09vUr8qf83gg/42/8PUw6Z/Uckz0LbEdqcO
AoDl/mq60TJC9OzBQ0fp6REU63QhwHmw+QcY4Y1+HqQp6D1AfpbCvshHqAJ+rMZb
gIhiLFbJPNzG3IMB77fAyGMWOiyxwUHZwqzkLoFXdCnLSLovgc3nVOLyGAqyYTMZ
KUwIUuNmEl9k07l+QfryWOUjvF62onnPgngLvRYRuQvkPv7wPZ5GwycG0lE/vWu1
OcqltOo76s/qF0I1SfEz42VKsJ47rpbw4yrihKNtYcbJfyxCE2tP6ZzACiRShuhW
HtJAwsI5tp25pSdS6ukkFtZVS96jvFZcrSILIKhu0mf4HBN/u4JqHpFeGSEmPiww
LY2K61jHvDWYU54Lrj02Bva/PXS8dhCKCJmUiG61RAIlu9V1PowwfRuGZ1sAP9NZ
sevyqFkcFsurC0N/Y/9sFZrlyr4sfikxN2jleAyRpxlPOZXuhWMTSbD1imqaq3yf
Dr6aHWQTI2ljCuiU54XF3Z7G+TRbzxHGIC0OfGElQnSK3XVuxJPm1xUrRYib3yaP
EPvP4wCy30s9hNfOAavZZxlZzXugG/Ed0o99R8W0WfZEKINfVFfhOhCH5FhV3oqU
83JCMz3qxyaEtxoEDQ4iGqKxWW+zUsNwsDesHDZm3ZsMa0DmDiHXTelilFWspiDC
0Qi5dJ62LinfNDiVhPQKoO8+lVLL5/O30XXsS3ENQHVTQXciOF+ZCyCa/1LSXmMc
aTLg2Fc3X6RtVbsPa9lbGn0qjLhZbHhs48G037FwwgweaqPBjIPBpGlaZJG/zeYi
3JwbphYeUVzXsWrFpowrl5mX3QAARfVy4Mt6aPUD3rdwiyTbUQJfV7I3IzvlA3R7
I3q7tY6UTujbaxR8+U/QlkpQjOSTzkUjyXTVu8u6tlm11WwExZfCeiRcZoJEiTeT
q6c/zQgf7s2LVWhhXoGbXVO9CT9/Q5Lmso7tmLRj9riHt8J0/ygfSDT7eroN/gpf
58k5UadnjQM/7sYFhr8VvNmcoIm9SgV/Ughn0skfxzqoAKXo6/NFT9oYg4LwqeWz
UfNRSDRwyW9yrESPC6SyjYs+qHtmQXYY8jkTCeMAqf3s5H873rczgZscVeWobWwn
RZOZ8uksVGbkJ/c814/dWUxJ09fSf/5lIhMnlo0138PA6VheC7JpjcY8U8FXGvDE
XFRsoJ/jEJtUzqXVUTF4CBEIOcfJ8h1UgO6pZl3m2waFtLS9VO3vg66uKTUlySVf
CagpqihnwO6Cg5fKECo7hVe7sF6Qe+mUL9MoYKt9m14N4CNkyn8x7Mo1xSHIE5Iu
PxAwobJVJ8668VLG/EmR6dQds+bBEipjjg/Yszba8oghv6XajDa6OGDwe5/Qf7Z8
pq2zxIWHXrKDH+zBpZ5ha1YjLU6DUoobkuMl6g6wNZ14hgPP/ioJbnSkwo6ZkXwI
TSggK/tTJRcuiGxDHIKaFzTuow6RLVW9t3sWDBdaQA6FQ31dEcQXksVH4yEEVLMn
oY3ABWOoEt4HrAMXsVgf5+YYNZldZiPVJxOxx2l2OVb3HT20DIdba/uy7f/DC1Zf
2rsqFyGx6tVgOEpm2T9UGemUkuMtUZgq2p8L3r2zrwEEEo8TTevAmswwKFJw0HPa
MMAmZ9RgmSGGGgPsv2D/YGGzP9asrnVFVMCeMqW8YJKrUgqi2fwPcFB2cBZO5ysZ
mFXT1vyoNAWcSi8r0mMfxemkFaM0WtOyhoLBXCncxyJz/1zSMz8a4dIgacIv4Won
s0Mkybt/UaYhcEcfZb+MsMD31ZsDqm4feRlbGFl9HoMdT4w54AwJIGJRtkg25va8
59B5AEJ2E70k9Pi/EgfhcOPZu+rEQ27QoTyx6/AB6pQLW5aIwbHkqXt9UhcDrbvC
35K2puFa8st/lKU6MNbp5ydtKSjBU0BCd8+1gKlpqlPwzhuMT7hP6SbkCs6n7Nwf
tZAL0X9c+GaMuH3Gs6voObIacLSeBHIyyhJVccw5fmqTlpHSCk57nEI9258n4i+u
+soi+LyCTwU7A91CAnjZMt2IY065oLju21INphHrg6z7kHsH6SDPp+gqFOHjHew1
7zHKfAe4i+F6+jR8mjk7MLZ0EIp0wfbx3SO38hNQXOAcWsqRCcn1oirJz1yvNYdO
1wmYls/i5ic2Asx6KhzZYTLubRyw2Xxx3YMy8dWm6BgH6eoO2oBIrS4FpFrw8P+M
botAMTJx+FNeVF2lH9jfL+qXuhf2xuLR+Pz5SaDELTV1KfrmqFEaEja2I6IxWHhm
SjwcY159WcaNTBL0URONbbH6Ak20I/OJBfGQwwIZfoRurhhTiPYQRkiJ1q35rYNw
22PXewOSCunktOkr4gXLmBmryXUkTVOI5kYtTlNMKIe86duIvrkvspVgKRF9wywh
elQh68T6YxJR5DRgeNq2sRL/HxAQ7YBc7pK4qnQkhYMlZS+7/GdlAsEsG+KxNFnX
gupUQVtmeLMrZnLLsyF9473eaMyzD7olaWdemzWe9OrqTL7bh0+xgTmWMoAPhA7t
0wjGseFMI7cZX9fJ8ZoULf/HYbrHvcisrcYsJURZy1nzHVM1YjZIWbVohTwJBBqm
kn9MCH2rjroYLzixXdadTlCpn9RyeCUJt3dqdIAGcsuZPxWlegugGNZCpTeVT9MP
cmMY1BUBJ8e8Tmyoei2ZWyPqSm1pKGTBcga8RHTG62vv9hTZN4D4OL06Oe+MiM3e
eX4prfCH2rQZ6kAwfoLEOENMHQqaDrd/yeocldzUIBX0Dk6tbHxa0keU0cetZMjk
BvoqEaHyM8QrxpBdRX4W7GGDZyXktKfsDuerpIGg6g+q4XaWrMlUgbPh4FdEA1vV
QQV9Rhthp1dTXqNub7h9s2Nh/0PNX/dfNpcATFmjjGNSILTUUEq+8aIJe5w5z7IA
DSrih7vGon9j1o9pcBzvgQlD7Pgu5EFi4sZCVQWqK6StU4CGssw+koRVvm4TqIXi
rrnSbiC3UDVg+n/OqYo6PMOskcHuf8CZr9t6mTmj3pNsAMTT+0h2ugFlYTvOYztM
Nk/z3tevOqv0+UVFoaV9hiN7fijPWd1INrol3nKm5kMCri6iVm0ZBLfDm8Me6/rW
An8V1n2DUxK7i6yWyyDXHe4LvrNWRPD/DYQy1u5hK12Vre9hYCdCy6+A9jk4l4qT
uSHwBzO6PrN8VX9YQcP/HlbgpPYDbjCNqNTCBwkII8CrnKJisnYniJ2aODvRuqEr
Netbg0eLB4Kj1LbF05qTLUnoh9ivY6rVUVntWU1WFPl9IswhB3gpbPpVO6fr997+
so3Jy5KAZNwKJPf4rAIyJ9KnUotxC5W5bkfCrSYByY0bITHC9v98TYdeEb0RU7HJ
rse+5/x/tEgeZXer1gn9h5cu0zggEZbzSXZz51wd5fbVX3qrERC24LzTVw13/usl
EvD4+Z/8cl0K/YyYir2gPLvFAB/gR2Kt44HQBHP1lSAN+8eHInO26GWWAwEbLRrM
lG+U5hZyql2bbw5/7YItjxNKW+tAhb05uZ7Y5ewR7kxEGlkWyO1dRT75rFiPAyeU
DyFpzf2eEv1qCF1a+IUFmwOzCTAGogaT1nkj9Ct5sLPNx9GPt7KcqWPWit3b4iM6
cGklJ61ftnudaxrWpGZdvJYNNqJCBu2D5t54jS5+p1rnqqH1RTOoLtoi2fohENUk
jvY56cj5UaRJ8SATy1idh9wfHcP0Gkhe6GZY2OLo8a6if0GIXoR1s5Zj88pq/r61
NS5XOFvVsGx1/1VR9GeoikX7JcpAIOB80/Vg/6s6muCYzVI8NHWNj29nI7jsV1Uo
77eDBHDQLT/smXFD7Z2kXDbh3T7mcVBatx4c+q4gz6Grl7lONglkSZI/F2wFxDdy
rCr08VUK08l0S37E+pn0x81NR38WN5n3xIev6UCq7pd3KLsb+4w4MIwGKIxH7RXR
nL6o5Q1/k/s4z0tdT8gZUvu00+qjUBt2SK7Dv2fLrR+ldaiJ1Lls4wNusc9FRINV
GYRU2rEhk4je9Z4xgCzRIlMYvS8HaXWrbrIU6XSYe2l4zTLEMzA+wio/NfBZM8IP
rfUkz2axxFsCn878LyQmu9Slpm7e0z5Pv60mzlpCnnvaEyjho15qxAfSWkziC0rx
aODYXGoQgxtUUof+u7kYMbzPuTbbjh4SB5ndpYMB8rdm9FVlNtPWef6uKaqADBVV
TsBfQ9oWQ3P6cXH0I3+A0RYDNe40HrpTyirBv/iDxSvSl6qLMOevzIM9ecGYrX7J
W7hti2yuGUvxxOaUtx/aJlBYlRp11XnGJE+s79CbGwXlUy7QmFx4+Ecll0ofTeXg
W/PAa2/ci5LlQKvsq5a8uyqcoG+R+nbe1QqZVlpXCKWEONl5udmDtTNe5B4aL+BR
RnGLA9C0+DNf/R7YZfLPZOX1YFSjtm13dCYOChHR9C7V3rWst3nEX7WKBbkMYKQN
g056MfhVxn9NtfrNF2YW3jsEXZZOM9ql6elRwL5MnNfvXNv06QkndsjQPDjaDpMn
BMcKCM0d90DbhauaeERR2bSbArNUsSgDZ7PCvKI3Rhu3pEzIDKH9nv/6he2nb+c0
YIiPhZzV7G6GbYSyM76lpfqnoyI0DgHgQE9kgxVY1h6MSdIx2InmSMss+X1RRJ3C
EdFNsk0uTdgaYk40fZAeVzmkM5YfVFQoApV7sD9SM2UB+80Sf5hJrObqDOx2Chpy
tZRCn2QUZ8dcE4tLOx1yD+QSSWeOFKnjL/1jg9veK9DPz+eP01EUm/6FmqsNptWv
EY4w9ibFEnawMYl9kLZzRuVtIhGZtQjDR2oCSe5WZbC4e9+ruvjdpccwbK8cEPEd
ZOD8fR7/q4EmpiWCrgF8dj/4gzz2XPDURwBnZ+JBJLvkOtbDMa+wNxzo6FpJRI91
4FSHMavdtgupJHlDHHRSWrfPV5ameh93TWS4qW+DIAGureBWn53OrkME+9XrgFAr
3oZ7CPVPUk9oFcTqmhHJfzOXviF6FLebIg3x3ymwqqDBsmVXDD/5zWtlYxJNxkjM
ZyMC3hvW0Hba8gxxIPKflQpz6fATBnxgp8LmiK6HJOxqcOP1J5Qg4xmweUFNp2oj
qynJ2vkBq8okiTg+FcOTrOIQMdvxrTSPIP30HySoEmf2eKGl4TCuiTAg0fF1UJBd
Dbi30XqwXCvtqA9bZxcTX9TyOh/ek3D41xzMqGss0RZkhlcFlb3nsm4TwbmSjbxx
fCqq68yLQ2prx/qPmZzUAJwSGSxStWvgmApzutfImvm3vBKGHslPRGUzK2qkS8Hn
R0H7wdcod4OZLD7IVt07Gz3KEKmMMJv35OcUMk/fkFI37Vb2/zivwaICcCBUIoGE
8inI7Vb5sh79JgN274uUUg+ldQoSXZBs8owrspOQcOEjxws88rTae0Tc0Ouu66Vx
WlhgdIqYywhPNKWL9KPuk2AnSFd39CyTj7QADxJTsYB2SF9JtjqaWCFVTtv6kVCZ
XLSNAOjN6NMtLMwugN2sJKZLXCAMWbbooSPSOuA/9MT5pbMdnyGcYljfDJ94iWyI
qR1FS0dzLK4LrimZhhFDTeKx5+aE0lhd8SjFutetO7ZPZ5Mnb5vSdACAhYJeDX0K
k5EJegANefflLfUHbeBHsMBDwjPpbcMsqZg3fZ2guOm3YE79/8pSNCb4M/GesVDc
x6uoHKN8qdFiJB9iQnTEDu1GYOKYUnvojkRm8g2ks3gEROr7sfV1B4KrNbCreRG6
n6kV8YnFaotWbMAlWLrdyusAZMBa2l5T+Ckg4hZpltpNohB/PlRMp/fXroouLWk7
zXiqeW0+6s/Lc83BmLhf7HoiDbYAFuVdgpr6K4osPwzg0HndvujphtDuhNy+7KiD
lkP7o5A7Ljd/cd/qeOYVvn+okDIgkS7gbtLoCVEKTDUJAkZuSPWJf+YPOLCxljMP
aYduJUCdUtFvsMQP/SWnA0tSobTXI5ueR2NHNoZBPkYku0bdat87/q02HdWsR+ki
2Ybkky6wPGFGjLJrhN6GMOkHKLBibxz7Y7i8fCL7EUACyUrTG6VY5ra4HvH2mxCE
ZaEtEWAfuASpLweZPpZfC5j12HHBPd12Q0L9a0to1+i0brOHfwJ8KQZOR567cGBF
X1NgScrxflK1htV7nnsi3UbPV1Y+4Pglh8ZXOMPGU4pVATCxaAN1mLBwjUsTEr88
UzeuAEiLaswU/T3wcdLAdCXuV7Wrpv2dMHE7K5vXePABjaSB+0wk/2AaLDzd/y21
FbqNk19swD1vTSr9krqWAO41ozZqyewNr/YCUGy5bHwCADWJLUh3frUsF7G+WDyp
xbloUZ11buNFnKbeJhnVYNrfVVDbnXftw2YCRWmhQ6HT4KpC6tTjPaggLLPrePRl
bU5eo07jgc0n6tl2Ai89s6LEyenY7MTHu/QXio+oLQgYnLhqsh1Ss5x8R9V5MuVQ
mIGZFfViFTMOeotaOEa9akZV5cWZ//D4kZnMkYEGeZtiubmcHdi3TDZptrhTbBol
11pffQ/v99FaR+gadZimo2dqnHMRAMt4U8urgDkBqIkWbFR/TanCpJnptyikjMih
41+JBRR58IUvlob4Rq9t+ft1hFzEiGZhbAxYTipKbXjP2eJVGXduCHbRmXne5ZNy
A1ajGm0ENba1QPfxg8D7BHoztuXAEww3iLznsGktKM0qys76p4WMHQrHE+99mAPD
oBxy9H5igrrqITS3jsrkQ5pTuOTfvsY5BUceTKo1jrpQtPWEer4N1kJRcafZhbJA
vxijr5Cxq+QBLprPIFE+8wNcyXJBeSA5UN/1BRdCFGAt/cw80FUM5EXv22WAVVVx
jjmtXfMhFGBodejH4dhaMdzOazN1jlGfBK4DP9N2/5EoacXPe2jgjLRnXLUAFQAQ
T8ON4g8aRL/i4awtY75JdKwwSEeUgV0JB09xkfjzF+HOixTLFaeGoJixqu3d5GQ6
xhofQ13OYHgEmtZW6/9hhR8J47ovhsJ/wJMDjP+j1tGi0tIqajdZYWJK8x8gRRzg
5Eb+fTv6yav+m4bb0SWEFiAKyy8zjgE/L7ITEVRysLAYDntrEbEzD8lyYP3ZEXPV
iG9iInZDC7j2AKdRFm6HczcoSOHdg6HK+B4jg373xVNJzsJKSC9qywqo5ZmfNRfB
9y7SbdJg36PZGL7kQNr4sLNRpqzAiC+PpyKaBwefsyu1iLMK9XAXhC0pmngM2fRi
51J0LCYqiUO5fFr+gfJHJD6zWvUbQ7vGHrvNK4Mh03cKTHJ8KluIeyjvD4jxgxiA
+4NZv7z/tm8dT/gRWF83rp55CWIOFO0bsdiGgKmBn2yF37yZC44ykxQ1LGhXvrJG
Sf7PK0HKTNGn+SGmWYHVKVUrwVwEM933jagWtH8XfYhCCGdaOYGG7oRf1Yd5EUNh
gOf4Cy/y42dwdAI2cq/pBod8rUpyImk9ihJTxDfU4nuwoWeYRJ4O4LO20kR8fTtk
Od2s/n0SQb7ogJcxpadOzbmD9aZOPn6fITFeBQuiX/JOk+P07aRbHPv0E61I0/FU
8d50ew3XBVWO5Fg4GJ3DSQSikTarfGyznqVavWUKVfGBwk00hGO4BStMI8HTXXcF
bL2ZkIslKYHxukBiAM6B1qb6nduwP8X7XEUZ00j1/e3PNuApCqCTRzNzYer9yaiC
HVe8DQHHLh8e1EsCkwv07uYzhKnweM20vmBBQf16Qrxuinq5tW5GOBPxlxK1NTZE
zdZrycc6FI2/ZbyaKIBwy7INLKMaHKa4Y9+9gelk/a9Qs8dvpHfJ4IgFpfD5CrPy
LwquNfzu8jS1ukmXGDunaeq62uoYyxFrLYO+dJYP+JQ95fmo9LIrGosIISZY8xrQ
8M6GmhD3ry+OOwUl/XTT13mlKkYhIBFWtyAmE9pFnIqcdCoS1airG47A2tx0qKPD
wtIH1ShqQl1LMvE4EZ6CfxIwUDkIo+CvlDkxGT0pD0TRi+pgJY2DW4enaVFZ0Y+4
UGGeVgyy/VdY8EWDVgNArEa4oj9tlX5TSNLgNwPTAxXG5FtZq05p8YHfmpeDa5TM
25Hh7a1iYKJ/sIvGJncaS9k4hQ9uRlCD7xipf4AhBzm479GHbW7PJlysgRz44+WO
ddUvo1q+TfY+72hCjVlYQoQ21ZJl1uGKqLL4C2AnRR5GGobsm+nmApSX7uLI1Jgh
l1Y6IAbhzGYWU4mm34OXVggn6YFwGY9lectVMNVIl8wPjVuTFopEcaTIbN50t9dm
xLitfOsXmqVINkduQ6FwBaDQESAI/2R4eqyXUHo8ERpbrMrYxbBBDs3CeDyls42e
DsMdSer5DbhzFSDmgQUPeXd73mZEBKGDPbxkrS3AkfikCrXz9jAcdwFiwNVUQFAI
7Fl2ogx6kX2lq0VVYzkXdCLSbJ7e2FmEv6IbM7+syXRSmgEBXeQqUuQ26CveCz7D
QM7/+LCem78Pewk0Ym/xZYG9NerFUBHMdMjVnf1/vof82kiTUk2jZXNWjHIutajU
qMywmNJlP3w37ptaRAUZuBNMYcSbf3rQIA2gM2x2RLgUuXVY9CXOfs7ZqMeu1VV9
IltHNF9wXwWAcX5gbtXtmsPaZsYK4rI+jsJkKt4epNXCHE/KJn0CGR1mZHhLlkRt
T+/2+HJtwPKy1WWXO67dBj2Y97lL5ySIlem10cq6iDFf47VRqkNZFBvqVN9QAvgS
Ezrr/n6uRMEbCWAu53v03TzLj6HJAZcKiNUFFHTtg72RGDhkY6yMSmRyxrkdL2cz
KKC5AoKWe7ZG4PJOvtYAo/aaW7ykxkyNZlfkYRUCfftEQfTbYAjXnG/SWfn8aVnx
hcWf7FIOWjm70oSDrnkfzUyRysCParknRq2DL2CI7RKwdRkb7H6Nj+HBk05JaSYS
/0/ZoSSuynLMWmX34tk0gCmyLMgmE8tDJ6dw8uscurd6vG/OtxwuVAVoslXZCFrh
xQoXhiBf7HoWCEvJR41QWw9rIPHycKob5lh/H4uW6lAlo9rAfpO8qZoP3cKwCnsp
RoSqv4kfaNlEI6h/Z5XdUMVexfwceU8KKWCvL91FMrwUkI8triV8DqRYy7imkSPF
aB667/FEv2n7debMkm4erIwiLHgAuybY3yq9ITpsJmUKqPYO3gTvTcfDlE5Kq5c7
Xv3esdrWEnLJOBmw+nqLngv6y5Ub7rGO2KB5Vk7Am+eBJrRBcQrW0n8ybzR6ofIC
gPPasOmlM+1Ij272CpdsKy/yTUqAAzCE33SdEgiJzzP/rrg7OTdzKyOg8qczw2qz
mv/nRD5FSq9saA5AdtgqWE0B4BX3fdSmZ7KFeGwxtHuMvWbH8Rhh9BUg+fxcaDBN
xFkFepc/vHxiXyPO74QEekuPw1mPCTTFzI2dQ9+M5HhEAsNt2Z6JHWkkPnZ5SvzN
N/IjpomFMaT/G9MiYVGY/xV4jVS+EeYSw/k1F0Kk/xfa7lXzRzdGtA8x5mMikU0S
TRjsS+iUncqDv/cppHtpyM+qfdXGPeLe0etYOjMoud0mixbfAvq0jC0z/yiMwJV4
m6o6/OTIqjJC8UeKb3SgHgr2VN3zKoMkw1ZPcrJ0hC446cIOKRupS1rHMIwD46Mp
9lKO/OP55E7Ct3DrLFHT/NN2DvMqmvaEhXSeYPE+Fg5wGrd4k7kEmQZC0mU7Yoy2
0zMaaz/3scFbX2xPI9gFHif/+pD8SySEs4iEFXZ727Qfyozx18RpV6lSZCHyfhzL
kdmfM03PIyC4jAVPI4578Q76UVI+2L3HWYEpYVXj8yoFALyCtA+LvsPlgSjsJJ+Z
TjbJmSwl76ycVb0eDbHwjrSiDxbtzBwR1yEHDfQhGscmIQMENi4Wc38dzv2rQRao
r/OyZekvFB8Oa0gkdJ/w5CtZwXz0nXxVhKSEJuEd25NdbjSnRP27AykSGq3L8oOk
AquWCu3/zfgK1OGKerWnzOcslK3ACQsBMEBQ6uvGACbkbrDMoLhN2ZZhcVb5o1W7
HXDm22naReNHWDIm4UQyNmiLuBIOG/i2IGSCqymbiV3UW2pa9oTIok9GOhl0Q7Mx
V/IiwefT2s9RmtayDJZ5/0SoTSp4nPMkqXELUjPI1YpC218ThOCso6346YFugNP0
0hqlkrbSEtVW8yZE1/wBZThAUqCV5+Bu3NdELtbUk3rXcmCEZDe7MJxsmg+aXZ6C
lOlvOW1AhmSljBAyQiQKMvz6k7lo2qXXJ7leBkSrV8oUPZpxP93CfHRLweth1DOR
P9rQiwAV8KLxDv517+4H6AguJFQAZ19sjK3R+l6or3mbT2l82HwAlxjvr+gg+vYF
nj3wTOXQOMptA8ZyMLdvtwcU/jcE5Y4h1O8e2dhIo0gXrFNznPY+pCGW7wOsPH/Z
qUHEPkwr6a9Lr9Nj1nIWfJWPHgIzjKt0muvB5eYJcWq8Umyc9UhFrfsd4U9emRXN
CkCbTwJIBdH9gVePyGNTynL/uC6mUlcPW8Nwka4OP9pKMapFBpXpOB4AE8xt2aF7
4TQIT606RXR2wxvCs2vbGvlPDDfzb+Zt6yif1apNxYTNRsdQmd4dWlubQHIN/M7f
Kc+6GpARcFuTI2p32chLMyB34EuM5tsDQwVY25mwCOPwP1ABIWmCFFv5xGlP0RZs
Qg6tM5FFCnZAl5txLrGLsRoWYKH618yaQJ3QahkUbljXm5tvc6WtZKVPS5jnmb4B
tecSXk6P3Kr9GKckw3NV+4eY04uKWnC6tMH1VdUxh/O6AMLFZvRvjtwKbDoADYDx
saPLxTLfV3gE+0poFc8f8FuspYRvmfO2UmeAY+YyQfEQKK3TNaqBbl1PVGK3nGrU
jbNLa79zWh0cGwEyH6VMPjmWYwXIp0mn5LQIxS+5t/4Yqk5Vqf61xWlhS67skx84
BpGRC1x76r+mEf9b/gVpUevF1kfj7zUiYWMcxHcvfdaAzX0jQ0Kcqwm38j5wu7Gu
KgcIDBKErrRCbDe1ASTsuUMreQID0vqHzcuYk+OEzqy5daYmqFdrVf+yI0kjsNaW
mMECa55JM7Ijb/fONAet0h5FJ5K9la7dpSZOlja+OpA0MYujR0cF/Fu7tgO3P8w4
POROGEdYZZ3kOLWfgDtF34qXwWuozurUFhg3UKif1fCkkNQuyWZzp1f9DY5sCJXt
ac65GwGww7NHfnyZcBw6dVZE1f+Xz89R0SHjJK15nzLWrBq3lAYjVltqXvlwNsd/
MmmqecLdHYg2lGxQnCxX6pJdUNRGLxk0YXiI/MSBKFNDDF1fRgtMY84J1ma5JFFI
nB8nRyE7h5z7NzzoDpFg90oXG7WIfUS2t/kNiHLJbM61oXbirbrjfkVhkC/PVVzK
V775of+10spoNBJQzjJAaDjwvC+W1xVUT2ij6sOEfyfNuKXtGgOhkmlHWHkPBJsK
wLyyfv6ebSerzrlRkwHXefEpBRPdBbQHDrH9U4lHEcuGybekpECvcrRXwcE/9/sG
eeJjFa+rlgJ5rW2fqL1/qRhgx72hdyB8/HiFrgTu/sj5l53fxWwZZw4uX7mLYWaU
QLt9Kiaho0/HOBYeMq4wqu3xgzZm0AfeQb6JGpfjJr8u/zZVxiomHtwZMccG+msA
/KXca3ENPwW4SEWanyUKmoAjupQxDz9aL8eQs09H+e9RWzJb35N7kBs40tjtuP67
oAHePKu8QZ89EUTK092MwVQFzP8fkLEjL0OPM4T2FVMTMhhrYCrURxKdJU7i4Npb
MQOiEMBCpUDnkR3qmH4bxRXKwlgJt9HgHo2ixn/F2LuiEom+wkshaeejVPFhMXrx
sQwKlZ3oIns0TzpNt47IzutSerxcONSDkT9mduicJqVl+qogAWVKUx7eMY/diMeT
QKSi3AJI6lb0t/b7Vf7vdd5W8lA0KXXmA5IA15MebMuLnsb/gcKQsVY9dsaAbAtn
feckQ+p4edmoeMpIZx5xfAJTMbCyoWPKliqlElCRM4CRts7pWS6cg/QN6NmuMeS7
iWzaCUEkqtccStnt/fRU3OGqZMtNBGukI8qmCDGDpCSLrSCT44BNKk0QSQ8x9kOa
hToSaVxGQGuF3OhASbeNH9pKSsWSsAYUucNHbzAtbhq+1wyKJplEBU15wId71ATE
nTZfcklymjnGW4lp2PwrXzu/YL7ck4rvN7mY11dBCS9ZTWLFaNV3m3PTiJzBblDO
w8fhkWPPcMMWDYR/d3tZGrYpstXzl9Jj0oj5kxfkGUN6sIap6GgOo8FwRjZ4eF3a
5p95EKsbhXXOcZgSCSJOsK9grIkG9bbbGpjEXvImwYChWK04Ce//RVUzH+URDyl6
hRrBDGY96tzSCDu3j08ZWa1YgHAyi8n6CG4vUEuqgHlaITkyaogKnN+6KjjR/UgV
lFXi7oz7B3+g/DkhiUGvTIxjvKD6v/JmG+dTiYncDo121xcu61nftSz8Ms6CI5At
MoCWgfPwU/TRyDM01AUnwM2vsUlGqQycVTVZAg+75+4wJXxHPvp/1FCsKG4KVCjY
i7SE5Uj+qaKfGxKK4TOQo1aaGat41nHPFe41pM6TEsx0hiYM0tXTin3iT2YiOahv
oMhurCl7yOlgZpAc9DXb6j/v5e46IIicPWSxIZXkjJ9Vb8MwAPwamvZpmQgCGjf+
19mHgVYERRHSozhpD6yNbWk4/tocaLK59DsxEqOc84RLqn4VplGvafWFP4mp/Rma
b8rjjI7JJEi/3uDEx5TDCqaAXoG6Ff/TVxv27/SffCQ=
//pragma protect end_data_block
//pragma protect digest_block
eaOoOtm9dk23zfCdDdU0AklbsiI=
//pragma protect end_digest_block
//pragma protect end_protected
