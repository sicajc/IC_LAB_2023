/*
++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
NYCU Institute of Electronic
2023 Autumn IC Design Laboratory 
Lab09: SystemVerilog Design and Verification 
File Name   : PATTERN.sv
Module Name : PATTERN
Release version : v1.0 (Release Date: Nov-2023)
Author : Jui-Huang Tsai (erictsai.10@nycu.edu.tw)
//   (C) Copyright Laboratory System Integration and Silicon Implementation
//   All Right Reserved
++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
*/

// `include "../00_TESTBED/pseudo_DRAM.sv"
`include "Usertype_BEV.sv"

program automatic PATTERN(input clk, INF.PATTERN inf);

`protected
73L>aD2SbQPO=>#0:UWgN:XU^-^<PJ5X0>dG27;)0&X[3+,OM6M+6)393V_(^U2W
T33a6@5U^2LV9S89<1M^e8O[QPVeXV>QXJY#C4K)NaQ;)LF<_1UOHFE;+#6XSB3(
V)Z).g\/,,UZ5NY-.&gT##.WJfC<;Z]&G4@&<[e:fFbe_Vg/.1g(R;[G:S)K-SJS
LMHQ+8DLCA.\C>+P:DGaMV.JB?XYRM/K-Cca-N\H;Y[e7+D;?]@:P<_\R1\NG8<G
09L6)R(VU[fNN8cc]^f,P^6@;eRRC#\HX2CQXPME6:8E_Q3Nac3UBGN=H1C5D]g3
\@.)^-^UJA5TZ(fF2aUfQ#Pe-T6W1L\MBW_J,>a\CaZ>+dAa?R=B=/]>F+6\Y9/e
5g5RRUd5cBPb=PKQD\)TfO<^HOW(@AKNX>_K0^LEE7)b)EE5\ZLZA-6,?]e_)^=0
+D^ecJ;c+JJ5JBYecW[\/5B#E7)2B<.O)R:N?fV4:4P4Y]9UQSJbZTJPGGR[g3Wd
GHQ90_A^cU7K-VCYgWVV9W)4;IGA+Ycf87[MTRcMX:Y,;TQ>)F7_<4UL<>506,(b
/Z7TV=35Q0ZQOcf]CLQ?-74K=f\L(Hgd<e4#852+X85KM0\2I)V5,Q0JA+-G7S+)
_g,ESMWMCSLDZO7??a?,@[-9PW&>aQZ7XK5OeE2<]6=]I.ZM<0^Gf5U56b:aUH?G
<cU0Og_S)P_[R5SQ(@#8#4@bB@?/7b>bD5T6b1c:PBXVD)ca,eXE]\bO0U__U500
P0I+B/3EbVLOR(E1,37K6Z/(5N@dM33L^@4+YW+>D2A\:(HO_]PVS;Ud)P866ALK
->E&BZUe5d+3eU52?:3P2Y(2M19EeC,?Ib]25+H8#-OPD#8=JDE\,8^J,>4@Q^W3
N/<5a7T17SYc:7;9e;K]6[F_J]e:\>@#ZbFZ^C:5@T[64M(?67fc<LS#XWP+HCX7
J,@UDSXdPf0DO,PJ@Z+<T=?0&c/=^8b[-bC8K<^YPXMKC\X1bVMbWbNg+Q.)JZWc
ee>d(62JR\g_c)E^#e[NAXR0_Z@#U>UfN74YXXUIO5WKAe60NBQ^cL]5J_Ye:-ce
;VADd)9ASZ/Rc?CCE?ZO:MB/eFEB8\gd]FR3^c&2X6XegEAL]X.K_TGFH>Q6217c
4X+=DJTeLR7K(EdY_]3];gS071+T_E8;1>(eF2e2:[P@S1N&5SR^EaYD,_8NNU/Q
101_8+PaJMbLS9a:9.=0X>3^A+\AT/AXdWNcDf5\8X@H&-ZQ8+;<gfZ3D^dNGg8.
&3([ZY4Ye-G#M^aAO4JDDO;.X7XRCDF(?1MD<A()[U89X)Kf6^BbHTBPSXHDOR/)
6b2g6Z5-57G79@>=fYC8.&SUd2([GV6(7IV?<W)c3:VFT0-J7^P.\d3;VKY8Y]<]
G-,QYg@W\@d+PE;I5OJCdbHQN<@0[@,JEB29-N@_Oac&?dGfN.eO?O;_0#_=fG<b
0MI]4da&G):R]86L:#AZ;86.&KRQ2Y80:^,B/>>4H6-d/H?e-G(_O3KQCDO1?&]@
^?I)A[Ob&XW9ad9:8Y^09@IMgF9g=&IG@J=3OT-^9S7O>#PgFUPb&[Q(R0<0:-;Q
GU6OTS&c,A_#T1YBg0@FH70-c_TQYY4.YX<IG>WcTV7FP\d@-E9>=T]VN+Q/ZB6?
2V84HLZT#<]T&LFS9&NDWP@NRKabR@QWUHY-F?IGV0G^PeH2Jf/Tgc)gB[<((A0b
]RC](,8,=^PY:U0JL\)F0]&2D,^V:KP([Ha?2ZNdM)fDMY1:Jc(,W,=?KO2JX>N1
G.B[S-;\_Z8<ZF<>=e].SD\GeS>-_)6WLgT\^I2[PX:8KbF>WeG7(3eL_K]Z+]UB
:d4e?aVME-6#]+]M#88(:eYED^K+WeJ4(1\U6+W0WY1L9,8eYE+,>Y&6bacSb;.f
7@eO22g3,@ZJIH)<eTX]KcN;A>SYX#_-6DQ7_L6V5K1Q:#_#YPE)SM#X,AO\:JKD
c6-S]/C>6(3:gEdV(H55L#I>;:TAO;[#a#NTEEV;+Y23:HEFc]ECH]O4AJTe;M>4
FW_Q^:_[=)<P@a<gDPe[fHSRW]+@aO?O[<#g5<\0ST1&E_T[Z;=;bcf1Hc^UH=EN
K9?U#(C@>B;638K<L.1IZB;(5cO#KWX,3.F[)>CTQRf51#=Q0>G;V(XZZ]a,VC_]
e]L0Ad_e[D\<CM:IK#-3-KNOD^<abV]\F]+9QbAaR75CB0:I431eA\P)YEZ=#H56
d#5]Ig10CQ;c[/DJ.&VQbYPUP2R<e6I_(9^PK@2.:ggL5D31.:>)MDdLAFfW+KgC
W:3d?fa_@_8L]2YODNS9aV>E?+R\UK0f7Y+<3=FYT=>LJT,8=^MaEH:US/#R+c&?
,1<(=b1;Y;C:g7E5A+.DKD7KXLCFDK+?C87?f_#:<G]ARb>0D8V;,?3-4I0)S5]F
E;<_Ra<\#Cf+ZebZQT#G8@a0[X^#B]H4G@?Q/gZADcK>E(1\cY=5NMY.S>,_ZNQR
ePZ^PF98#2)A5W[6ZPD,7<T[I_A9(@HOUK4#.N:/<[?G:eSP?(RELgJMf.N12+YM
E?30LSK=)g/NUJ?^U,KHJ&cX3Z-\H3a5L_W,KRBF2)_/WQ()4H)Pc9F5G[0(->cS
d9D8XV/XS6D7&+AHaUZ,R-I_90N^GY3&QLM.>OeZLR->Z4OG^gW06[BWK7M]a:&b
THLD^d?SF@6GS&]K=4d<<#aQXa)):Y#/)TKHKffg8]-)b-,H-.>J5(I6YIeD[3R:
aIAYeJ5DNFMG[C:LRW[#Bb2JPY51.C9B_c/V.PIJ0G(fZ,5<R<?T/(YP<,9NM7P^
Ncc.;CgSPP&W3#93Ha_b5NgC9gIO/JP6Y@(KS@>30.MZMP;VS](>@/-+Z4,gH9[N
J&=ef_]fDaU[]LJU^)c8W?CcT@B9?MXPJ1U8OVI[YE(1NVR/[VPY0,?GKWX+GRV_
)5IR-KgW?aRUQ7C\4#bX-IP=233a.FBYG(:2eF_4?.IFO.b)71R5=/DbWT#aNc^2
II-#H.XQX2ELJIae&be.1KcMY/GSC.DNY[Y?7JSR+f71=YKT?S8A:7NN,[;^;@/G
LO-UdL]DObOa71bBBeNJ_N0PG/9_VW?&Q\,Bd)4[09(_VNXQ1?^,SfSPFb_6ZU<E
a[_IbP/W(I;VJ(?)>b]N28R1b=ecOF4?9IR\gF0bIWY[W^@M>ZM/[O1^KT(Rbab?
,a,\JJ[MH#Y:[f.Y<ZIN@:7d8B(/Gc+_U26FDS6>I/7XD^0H7#dU#<IUET7(LR?<
@BR?a79O_/^EMR/F7HOCXbZ&Y^O[bfK.9:M#J2D#L<^>7K1F<NV&DAOFT<OWdd[M
^1TeJ#+BZ-=;:TEPK.?TIRX>_5MM]Of>D7]-+4d;F,Q3/^>PEM>2=KTA+<YE/=?K
7]SM_;RU_(UJ)7<;L7/fMKUB7fXd;7@NRO_,9D?,)[3?>_<[d#KU?VPU3S_W_=Uf
@\^D(U#4NJ;(PV?)&HND^LUA8]?B[X]XCf??Z0B<bALgQU:RLdgb>,@7B8Sb_+)8
+6RFF2dOA64-4EWKBTZEY#P/Aa8V;6H(1O.];JdgQb24)?]WV+GN=?R5:URVKJd)
Q-^Se@;3JSQ^]a15-+-LFWU8FdHaf.8;M-B_BL0H6e#(ZJ;F^U5,a1Z9<T7YdNdb
2I;=>3[]agU7_M+fOKS9^@]VL7VE;O?71\R@ZE1VdT19KRK(/f[BAI@U;199XX/C
552f=LQ69GXC_1aU,7FQeS^eXWMbX\&+d,fP^JG,B)QRJ:55C7Kc+@V(d&-LQN\O
Fg7-2Ke^AD];aLTRZeJLU;K1R-EZb8R&;5W=):<Y6MOI]K]W\2M\L_@R4FG,&M^?
/gPH^T]O9UX&5XV:&>S#?28>K\^)R,J&dZA\<fELgB3DggE0^AM?#2JC,PJI.?=D
g0\RHPgL<f\3)aC0T,VWV&6^(9NO@g\bF<O:5FW(2I6:.\.Sde<;\E2LN,R0B@+D
B,_;IR+8>aE]4EFI0eaG,8W:Rb7YE<R0=YH&<QK4,9.+.c7PaP9Q00HKI4=(VT@S
EMH1[[T8Q7+.0<#A9<d=V;KX>@f\A-#4ZQ9/MDC&:1,0Q3P;.gCbO?Ga#-ae&(f7
U(S32T;]>^K[GSOWWJURLL7?;GPT(XE)Ig=62L##74WHO8dF)UPNb#TU)fVcSA.g
/EWO8D&:?fMAOW0EDK#I1XJI\:J:fU\VO[8Cfecg>ADEJD@<B74DDG#==4OERZ4)
&>U<BNGCNcOZ2g5?e:?[R5)7;#_7=LZ@HT,bYCbI&[(,5R4f;:)1(U#?MgTH-SX-
IC<L7_3L2&J.J5TaIB\?8@O\NZ,@:&>eB0XL385:8FRMa/;D.L;:eGcC3SaaG0&I
S<SZ4dWgSfM:;J_=@>:H/0cCVAE1=&?#>5Q#B9+&ZFBC1KUB6G2B[]J_T2)@_5MY
5_:/:Y7aY]>:8,\G(S]?d(N:g7(V,D0=&98LXO-J/)@V&)#81&NbI:&64DTf0TT3
U):ONGN(d5aU-R4IWfKO&R+II,VC.9RJAKRf1H=FN1<7dD-[-&G&97eVg\/-V)<E
2D9<9[Q5A_.Oc_KF([7HPM(0OVE#UKb+d(Eb21YT_Z9<F_3A9[P>.5,=E+?eJJd0
L0&M926V?XfU\Rg;AB,LcgZ:eLJ_S=ZXLY\\X<ZFH?0V@U(b5>Z\/N:(>2cN#bQO
CZcYIZ-0E98+cc[46C?E+d9L^@Q(M=5S4USa5_.UQ=4gagCZXW4_O/fCQE0d4J1L
+K=+?:45E;=+RC,@_3.AGcJ]bd+150X(ZIc+EdXJ-Fd-=I3N:H;\aB2-W8RKT1N9
B=H11R)?NY6&7TIX].5UOd@5\5+-+@T/(X_\Q7II#//T+eag1[a>e[NC)2-]QfQV
?b8@ALK0/:SK-U]\L?NHS5]a(>>#]45S#ZH9>@1Wc)9>@,B^g<F^fKa)&RSAN+-#
H1)@S;OJ^G\28),.6acO_Hf4.>V_H1MHV[JcW(;dWdRb6(GgPX+QJJU:)F.:^\9;
;]1#cR-L9-(O6C4NK1B:F>20OD?^E]]g>;OTT&;T2T+Mc^^T?^MOT5DM,W;:YL^D
4&,2/:&V=OC<^D?#aU=FZ]F7Va6-XR(?Fb/C)&PJ6[W8KVF&bWb&XIKCYLL)G(:,
9@7M=+7&ZO#R?SDY#a@>\XfG1T2CYcL1G+W.=XL04:>_FA,fH2FV?(e;J]/H>HZW
R80HD:(H:3O.c[O;H6UGNgZ>KB.MNP8W>17(bK5R02A1+WJ<=CO?]8FJ,T41_HK4
W+Z83H0D]48+9>(O]:I:XVda@4?)K98+]E_LEECBd#Y)[1)?fW]+]TO?8g;RHW?>
^9fU@Lf;DSS3baZ1FI-a9FMW<BWBAe/_-ITK==ID;+VI66(Q5.?<LABf8cMCEJJ:
@@QTFf[?5;GO2Ib](E,+;Vd&d>9_^6)G,Sd-GJAW@^1X1-6;FDR7)+PGb;Uf@YEL
^4fL55].XfG8ISU##FD1C=A.Ia\OL)#:DcU0DUL_<1RUA3?C+e]P4N:1^=+KR]KD
X_W<^.XQJ<T\3[f55=H<3gF,a-[-^)KJL8JeM4_?eC.@D=RPDK>Z3I,WA#fEF&XE
CDUB=3>.MaT<eI<4a#abW]2IacB[#Y@BVgIB]9gL.R71,4)\._0FaEZ6\\@:,E3Q
>^?-3;]21WD2:DH5+?PCMV)P:S]Naa41c=I):Aa\P<>gM<P^>2fI(49g/ZSbaaXJ
;<.\[G&(aG:+M(J/J3SBHYe+J3FRPYANXgX/L2U,AHK<TB?SY7U]9f\05>+1C4Q1
+3PZB(Te0Y-MSN7E\\)aLHcXVD^V4Od1@/bfK_Q9G9a2?7?SCT945QOLVHb?bIE<
_0C#X&93B>9ITQ+SRC[]F=Q__:8).<U]9a@JQgKT54MQV^3QGH1-8T<Dg[[Ue\<G
60&c/QT@5:gX+L:gV#)&Ka+,-B1R+1(I.U4A3Ga7QVaIe4D2LBS9)eMVYUMD>(7C
DA\W/^EK9+U.N>QVZ7^d,:<J[0O#4BPA^5P9<[64d,S7P55;:-?#VUdO.<6Gf2HT
3P+^E2@ZD72bORAd-/e-8S9B7.PS71Q+S_Z/B-T]XNf0Y#&2XQ&7SPa9]&?X39NJ
<QC[E^b;FT3X;WFg6O3.2P7V4]?S6&9)#+ZO1_UMT-=?GEOEFGFS]Eb&-J5SY+b+
#;#DI7aF^-Y518]#TDIX[I3I3:I20IG8=AOA<^[2,0cPH2Da3D7MV78S>K?&&9\a
<fJS1R2ZMN#g&Q&?TIBU:a/TA\TQUa2dMVdd+FAeU6Md=/#)@SUWXYXf)J=1[N18
-?())f\.Y;LJ65,dOP&^aB,@5KF7T#=8HNIc?a5KX2:T;g)/CUMF_S-XM^WL<23V
S^c0_\X\JT22XY]4NXN\c-[Hc[3=36LQg?9_0I+,(.O,I4Y<M=bX:3K-37Ka<F\d
e=A]U,>&SI2=[TT#&1>8P^.P^?\4-5?HV1afBC[N,U@-4)Y,/[a4]D/1EG.P_H]e
2:>]V);#V4f>UG9[dQdA.a#7cX.\38#C:8:2#>S@W<+.Ca8>_b-I&9(a4\&-T/;E
7^ACT1EDdRTEGK8JC.ZJG<=CgPM/TQ6^aY;:#KF6XS_RgVT+ESS;eD,ZEe9R?#E;
b40;9G6540I8OHN[J4\T,40Zff5^UA&?aP+^)[4cM5-JJ))@3b8&O^aT/X4&[d2#
70-U]MB\[2(cSISeWHAU.P_1#=\_Y6CB+?DC2,==P&f:eP<SX6NUaf)[Y2/,DN19
T)9HCCf:aW,e2@fPGF1UOF(b(gPD5+8,W?3<:b6_8dg>:GGMKIbDEg=YA:d6c4W4
YXK/V6[bG8(2cZ.>N,BK9,I7_]\AQd0>]_]TN?6=Z1ERE#?g.eZ=-DUcV2D^0,b/
g.KQdIEYcUb_B(L:9B0[TLKC&OCJ3^NT9=<@4B?V)3fTP?)X2/)c.gaQZ0</Z@)5
#9F/<8;L_,Y/.0aC-\DINTaR+9H26G?<(&,9b:^;3P(?DTGA5:RJ\73aA8f^^gR;
0R\3MR589VANHD,3L7BBN1<1&CID@A]HZ30W&-c@c+dHfT&:bGXV8]#SQP[V-#QZ
]NCYbUCEFDU:B8.EM2?eA[>Rc0I6LY:.<1F6:F-J+RS+R;c-1DQCFRO<DYH=9/SO
,DUfK6;95W;GC0>R:13cYK/???f<U?.:NOP2X],A<=OM^fHSeTE6+DaQd\2ZbFb6
bg9/g9W;[&V_&ce[[f;<g5C+[::3fAXJc.]DO@^bI5b](M1IN?KU)35XHRbd)5B;
F--G^@:?-1BZU5N#d.HFA\6.Jb/>=H<\T)0bNgg>:?>Y4CR6TgA\Q1O&?:7UTe[F
\Y2-,Y:8<b=+R\20g<E;Wg_aNfbH@R6BMPD43=9JN3#<W8RUGGBZ5)2#\dY?MXC-
_<WBTL,9,MZ=N.36YNc;.D2)5\01CRZ<PbN\@0<P?\HeQ0Ne_5M>O^7YK@3UB^+9
V_@6;HZ@<4TP)<-F87S3+c[B9<>)5U<De/+SIdd2AZ#6RTg<//#^OT^(JQO70,_)
]cVQBA_HRT().7^//aC>Of9&f=(1N,#6[H/G9TgI+]8^c<e8/(S/CBIAUU1-_X_&
>6FKRWNT2ffU@?>f..L;MAegFb5&4Z?8GF47BD]O9L35+1VdA-LKf]@U(^D4LJV7
(Uc/e^E5<P?+9P+W2)1#=3>PVJ9f2,?]=BH>\VTI2H\9)2YSgUUf;g=?81.XBagb
bM<Vg&M/MR.[T#>03N#6=M>[(N^T4/I&IHX5D/R/TI><TD1_+]c4KW)>?\B?[bUA
<AKEd3A;?B[H&R#J[IB@G_A2-Y]<YJ(;QI3(D+.F-7BH\d&JA)#5N?8))E4^E;M(
7L?2A;+1G=:\_5Ta(?f;N9d.C1HDST><]==c=]#K^(CW:)2UWQgM^(&;L/PGF^[Q
;O0.F#GXc07>H=A54F?5Afg)fZ1=^_f1@ISKM;J2#]>R-4aSAJ0RGU?4X_Z)\dgg
S5PBdF;e;O<P]#>3_S[KGRT(1QSTg>:(:=F/(\Rcc8DeBUaFI?BXcO&X82A062N0
JFD=X??.3=WJ;^H[ZW1J[^eaN;EFVX3JARNBCM-@=0->U(<VeASFVF,_E,2J52U#
-8UB6@.gDMd(:SDJ;U6.OR4<a+@6O+4XXMA0?P1IA:;4=gC3>S+5KC=YII,gT8\d
]9UDgE/1?[>VCgMA+?/G8\4P7M85A@ONS_;[I^@VJA;YCPdJQ7R4?P>.[;->YL@f
37fIQbF.]B]33HVKB<gcb-(XLGWB.S&/(BTY.=?a(EYa>>M>Qc7H>JKH&H;8B1e3
_L67#<L[&8X)Q1CC/9I6/^gA2V5e;Z0J+<K^OUeI(_.JT]gfODPUNH+gT#@CE8EJ
N+)4/>?Q0He(,fb#f;QG[0BB3-VR#P1HR>C\#PMfP/aRQ&[+@F/>]+CSaf1;9)-f
^<Y1^^(CD#Of7c/HRUMJ2?6\.-@g-Oc+O4+E16N04O.fV5L-]E?IMLOJcR&WA^LN
BM3>[Dd90<3c2JG^3bL.22Y>0U88UJE6/@#66H6fIPPW_Sf2Y;;9,P[USY.SCZXG
K.?HT#)Z-9>;G6DK(g#54O_1K0>^-?XS.0W=P__Ac^]=:a\Y=JOdBPU7aUdGEN,4
#3EL6<PU>+RSZ@PZ]D>#^2DAg)e>YM>\6C^4]+H_R3\:aXCL)4W3N,-.gQ,)VM>.
RYQa)cM2/97:[+PTU=6>0QF)gcZ)ZV)8(gO([]KJ/eO.H.KA#g^E)c>&5H9fHV?_
4]R&E?]:Jd[FbS00_Fe,9/-9]=GCR/+eAe@SKZ61>AP4+?WEdPB1YMK+9T&2#cTb
\4c>+cUPJ9_N99S/:^;1G5#V=]M>K@g5\KS?OaF]7FHUQ),2LQeEG[PQeX2KV,dH
T+edXHUS0CY^YG#2gVBbF^2-LB=eRFMLDX,[<G[dU-3XTKO1R2.<^3#(ZH-+AM8L
U<94IF:g4bF^XBR)gZK\=FSWI9AA84J5SfLYKHWUTICFRd?SZC._Wa-5de0a?7.P
=P&7a>(1fV+0FY]Z4G8<&U:5=cA7DGH+N42(M^KQ0N-+>UNfeKC<2d>a9=N#^_Ub
QR(eRT@6SLeH6M[6?IR]=eC19Q52fbOZYNA)2ZWeA6-,RT?Ue+f#\389U9?>fH+[
QHQc:SGBMQM4XGI[=UaU=)@8__AaW4Q&aB5O=Sf&U.g1HQ4+LbBBVF6b)cf(&Vd7
&:A:db7Xf-e:?,Q))/.88(ZFSG4N\U.aLU^].68?EOa?WId.42\\?g\;Lc?d&fbC
)0VgCU&e(XJ:SNU?e-N>-/^K9@KZ_gfWU/IC8X:XONS[[W7MJ(B[#&EH]7Lc=Va\
W^-fC.:d_DBUYQ6MdLW_Ld9-EV5I7(VgB+K=&S^>^#f[;cFM/X0PEdaL&bP5O,B6
RS:NeH6+cS>P?gVN>D1V?X=&B-R[fVJd[?6#Kg9O;:W:+U_@)Kc,dOf?FQM0)@E>
.dfBFBe3[PW.?:]]CX])Q9b99/P/7L_Ed>TCgIe7,@ce#=Q\f-TUHP.(X15-T5G=
N_&#,<\a1YO-D/O5,1MA?,X0II</Ab=Q.>[#9+DH:GC].ES_.&/)6]/+,;9#T1,>
a8RL)-J?[;\1502dD0A]+X/\6N\gFD[_Ye/J2DAE)g/:2dMb]FE[R6_aIH[S+<[N
/aUJ-aF@WL_6&NeNGg?[a>fK/TOU2KOJ8NgOI_eC3Q#Y&(M#9SfD=?)-5]5YB.Ma
AVN9?V#gA+FI6;eOI-:E2\&P&R0d@eK0B2]40C^BNVQC@&49DQ,a>&:VV@U6K#gY
M1_S-V+/>2+0P9WX07<^#1>bD;XX?g5/X7]^_VS-3BP93_#d>>W=DA.-f/X[CEYH
X1/7J1(@BN<[9+MfD.0\Mc/2/N,DZC)eYeJWMM])ZU]([HP;G+TRb</a[+VG85P?
&BB;0ZW@d6NRc2DMJM9,Y-e_13R/c0^N[@3?KH+7/MFGI9H-^W4Rg7.KZ\688IU]
9;AMdSb=B7e/He[d7_0#TMA+.bVC(25(_,5V-:9]&Sc<[;8dQ#=+>@Q_V\PVZAXX
PJO=U]S(.4O.H]DcAR#+/dc+9D#e6[:0U)IJDP]>G>fDP#JfQMbA8:U9_4=/W1?X
[aYB+4-T&a^]8AF4Q263,:gU[3<O84>a0YQa0.f3_g;7O2M1T+c:&FH8/>?b,V45
#Fe0QFeNL]4Y;,,L2J-=^FeaS:,Q()_SQQORUc2VM5J-EggX8)g3<FfgQ;J?6\8:
F2:O/F#S2KM=3&5H@@A2NJ7Gd,8U[>ZeYA(WDbd@LNH=b&2VN0e7CW+K>;/&YZ_N
g(:gIH6[YJY=c2\,1M)OH,g@@+.U=^5.\1/F+STW4e)G0D+NeD)_J([e+<M&;\3b
I)FaVCLYFYeLf(PTF<CeVIJ4UMOZG1FCCZR^J0C\eGV5C]8R8(UY\a1.C3Y^.VC(
J8DP_MRH27D+.T_?RJ6FS8HR,G^5R[,I1EM3[(]TH0Xf-Z@S,&C7<dJJ@,6-E-6R
a8U@:NOePAdL5^[KKCMKeUX)-,A12P-Q+_AK#cdD]BX0#&\Z?_M9OXAB3eHbM.PC
LAHFJ-(&_If^c8/PNb[EeXYI#^W-G6B0ON_+E[T9G&-.)M1/O#]B=]cK[W8V<[V4
T;(bIM=KB(/XT&AdKbG<:<,1Z#CYH1@SP[AJPKBH]?Rc3d\d61LLNMEMY_):JR8a
S>[51Q\]LITg:WI>OeO&964/[C8g,f[K@[0GK_E)D8V__8bW4VS2W66THSQASGRg
I.#_F@d<Q?4OOeBEFV=)=Z7&)0&G9b#V9R)+=33L,HH:(KR?_=QA<_DXa6-^<_[=
;LeE2-X<E6MQJ)SOU44@4>(2(U8_1=P-_Ug+eN@9&/?b^Tf/GXaJK@MN_<)9D]-g
:@-gSY]@+?SM\cKg];KAaM+Jc8UE8[P(TU0=^I@=F0JM[HNE0K#N[XSKfGP?AIM6
6^85<AB41,ZRJZ#.-U]RMBH@=RC5,c54@c7X]I1SE]_I^2?=H75;Y#C9<>JJ&)KG
T;I<>-)G&gC?Kb/;/&Y[D[&3E4?eQ7RH,&c.c/b9?]]O18<I]5LDHb\B[\C[SV&T
Z\7-2cIFe=c6:UL47FUcS(PMYP1:,Y05g:GTEN.&=GOH-B3E8T)gG2KWfHP5M12-
6/T[=MIT#G8PfJ9YX:E9fBDV=]8ZT(cZ)-abe-Wf@@1Y_B?&WF8M99HN,1cF@9A=
TA)cB@3UA)UN85PT_\ERI/.MQECTb:.E@3.Z1b..6R6L0QH&H@/@c=ZgSOb4QY,O
+N]B+P2eEe.gL<9T5&TWD/6L\KT+7W=9SdWPJMU?:NbUMR_J]/]9fE7FV];F/7cD
3UTAd7CVXF1&V<fBXcH\^O=>RZ=,XI-<1T6b=BW)Q#-3#R[WC+P)Z@X#QZcg&eVP
,d,IP00GXCIeg=bO>T.[<AHJMTa(EL-Y@;HW>GbO45326L>@I)C1MYLB.IV12ZZd
0+6#[1ZNM:f1725CG2Je2+GR@CP:UV/9:a-789ZFb\bY3G^cJ]12>Z-ZP][IV1NW
C_,WZ^U-G]+97Y:1B=3CKH@@A2Z/S=TS?@H/O@TJ[Hf)-g0-bDDZ>Ie&>8J4=bL\
/UbYB#+D/GX)a3;BAH<LcI7/R-Z4;d6MC7)VC^0ZQ(G=,;fW]2YV.W20+eD<;>Y,
A=W?6:8c9CG7f.C42TM.POLA4-IZACf?WO]P8)ccB>4PV.BVa1&b)BZXR.4M+Z-;
9+):50>P903FM>/V<8JHZOAUbDIF-Z/+3(DB]&Z?A?@[N_+(EU7=Oc5E3#gSN.S]
+,+=G=a8^4;#+4&):OQ\JEQ58AQ4XTM<)X3@Q&W@=,0OD@)(PIf/fe7RB/dP>bL(
0;19K?=WT<3A7R[G:dB4IH61N][T2J@KP5>-3E2?U\XgVCcN24+([fGBLIY=;[P=
5GdPd.0Y0F6EY6J1a7U,>]5,U.MILS)D/<FYR?\5\=ZPc0P#MZ8PXO-R,-J?PMS@
cM:cN1B-1N=Mf=:Ud,dFC67&1GI+>KeI(L_[\>5NS-U7Te1([;A/5ef:R53_S.O+
6#W&eAZ#JR<Ga=J/<(OT-<RK@8<>(HgX=dg.=B[,C)CKC(JcQRf^b4aGQXcA[SJC
TI@BM3?26M,2@9+,^4M10:,G)2b(54VWV>]a6NW0.=e)6;T1Y,a7#IB.QecC8#G@
V2&3BW5/:agc#PE(HA]6,K1]P(B@1G]e5&V,38^3R.eY3<I0;GB[(T91HO(VeV>;
3BY,K+(Y^V.<(\^3bY_,M.MS?fddbU-9b:;ZPbaG]X]J]/UL9DKXM\?<]W]Rf2]0
+Q?WWKV+X>1Zf;P=/E@E^&)Mf5XKg?AJg(O1,6M9QLDYK^.HECE^UP&B?[N+VNL1
L=aG,M&eg4ARN=JOJ9eJG\9Z3<6d]a.;CEIWB2JBR(0LFCC[8D^W+LL?L0N)#6LN
WF:=?TD[6RAAEa78X=>2--M(UH[&#K<PG,A)<>+(E\?)S:K4.PafXHd;56,_9R\(
5fY\=7Z9@ZeI(VJR&4gD582MWe.VMJYN-T)V<Tb^(/IN.AIU,#6.eZ6/37DY0G@+
\/RZUOg,(6(]CW9<3eUe,TYc(NK3AO1?62)5&Nb89^/A)+,NZ5d5eGB\O[Z9ZQ2W
+SD5\0C8LSP&K/.U=Q8f+7g;YW>7UT/)J>I2H6K:ae2OZWW][4Q9HU@ZT=TUbZM-
K/dDFQ<DeI:E<g@JL<U\2\P@I)Yf;1320(Fd>K97F-,A.ZeF,\CMg8IB^2R;,I+I
PS35P2O@\5E_E01LdX;ZCXZ.ZQAJKLG)b)_K7[2DS94PQ;#EMY2H_;Z)5Ma:I9]f
dR:789J,G99D6_.KBX^B07a#H_#D0=64+J4#@&PDb=#O//58A^NR4GKB,@..\1::
S:35:5>+gMCXQ_VMfTX9aF5a.4VZ[;0-#>&]]3@122E5_KbJEWG5?IR\4;3ZBI6C
I0>/BXV>T&3&UZ0PR41&882W+5C5Ke#K,+N-YEO#[T-B../TCFf^>&8BF;EF?K?=
e7/Q<JAZ2<\RMQ#Z66YIb1EFQSURRBdFL-AfIV:Lc:d&VI;(N_cSMN@7aTeed&VJ
VA.N&O=f918/TdS]eTS2AfcgIA0+RR6NOF;O<F>C1<7&5M^#5<T#;Y-6b7_>XRa4
daD0^Q2+VK2V7A0:9TbN=]^Mg^bIQQ=F?I6UVd:RN?#:@]G=</.([4D?YKMCG)C#
&TS87\3K1DBM)B>LLJJM8b#3,J8>&E;K8e=KdS5E=\0e\P;Ze[&_2F,MRR/Y(ae3
AC.P,2.bK,OIE1g.9Q)+K6YFe>?f_K:7f->3WSB8_FWFUKTIE#^IX3:^VUVa-c7Y
e-KB/=+B-aG@9URT8VQ_V2G?Bb_9O]YW3VPG5Lg8.N2K8T(9#(5N\#QS;AKAeFYH
V/JU_B[I6C.^\aJ\^V8Q1aF5DM[-5(aI/W3;Je^[DSU;K;U5(A\(R?P=I:5,gQ]0
F[M#GY2N-C\KM/WF@Q5+8/PfDdT#-.^=[R39)+_/ZS6=>\U36NZ;G-?/XJJ)EOJ]
7/2aIage?0M^7OZ94cG2I:(,PH65N,8S4=1XbG_R&0;=X21#6<K?K4d[ANINP_e_
eQT9aBfR8QQ?C<TY8f>?PG22)H8BBJYVF[+#WZ1EcWNC3cES_>;T[I^<<e/RA1Se
2dRQV-TOSK3<C;2T74-ND/C@H9Zf&Z4Kb^&U2Z\d\F8/0A?YZPc;+1>&/Eb)(B&R
;):B&c3GKL<F[Qe<4aLf9b>YX6I=C>\PGfYOeAN9@bfJI[]b;0+=W=a;4,(>GVb,
RDg:OS9DKMP/eVUYLOX=__\)4e497C7(6faagCCO/5=-BCgX63dLIRY9.=I5g^U_
.@f-(Q07TAX\(W=<>F1<2g7\P;RZNO=&@:,).?P#9,-6Zf1W/[8>H#Q9-Cf/9,VC
K0K2dQ<cXBDO@@+\TDL.]Ng)1?eV2H08\0JZ;>VR>EPXB[c@#9bG[HVMA>#8=R(T
<M[^IgVMP+M>KJG_^7O6#QeFCbg2XHHE56f9N&#=KK>0V\Le[HKZC46ZN.^?TF<(
a6.Z)8c<PI@>^\AON,L.,O,_8K0aH\Y)6cU1053YWf5)e;P=7e0;+F4d0g.E8H,0
[b&/>GZ7VJb4/4g>IBTY:.d;78WMJM5dJBHTR+e<&7&11IR<@]b)X2T[V[);0DR^
78D46:bW75L[XEB1;GNDbMH9<9@e>I#6TPe&7DUX-c+[322d6^Vc@BX2K1HA&#9D
3caDJY<B,dR14=1.+.fKe>-KN(>;K3^-Xf.SM1a^#P@.4RG.8d;Mf/?BcSK4aZ,)
BO,Tb5A2d^FWEcgJI0C;8I)EbdG>J1_EF#1QMQ5/ZMJ@L1@e,AL8NRJ2AG<C[dWY
JCP9f6g7J[RS]>^1d>1N+^<f#>bI386H0VU^;@G,]-V7(D(O&JI.U#WI]]UUU?/8
6QACEd2b_(ab=9.@Td-SZE0HK2).?EX9#^>-;F/;7?(A[1<Ug,3cVF/G9IR3?aZa
7IGL+eYc0NYS9+I52,aL+T.)QdDd[C40:V(87@GWM9/:.9bRH>HJPV5_6JUHS-g4
RPH1>,Zac]ZLD_ZAfVM5F6@FP+N3=XI9XF2]RH/HT_V7E.73DE?&=d746^D^T/YL
(,&TBJcHg&2KWD.7E)7:^b</\:[&WCA[6:bDN133X&UYNc^@E/N);dOD]c2PT:20
+KBFb.:b;J7L[,H(H\B@A,YM+LZ3aWA_PI[R<I+-CP6-da?NSUb,Y\FZ9D/Y/bAO
S1>1O@L9I1B@NZ&e19e^.8CVP_0_&eKZNIDb=YXK1:-GS^7<>L51-JZ9MTU:TNd/
I_b\b-S59U+e50(\bU#dgE0+(B5c^07_e5a34def/@LH9YLb5IWZ&@+EKH+1VeH/
H?(E^^5d6\d^;(fT_LNC6]I=UQeTC.V1WP/?OZGM1]BaX9cQ=>/e+Lg;#,^WU9Z<
f3UNI]16-f1-gV#8UG46@JVH?DZ<HOVG6I^Q3)+OH3L/4cS6)^6>@)CX@^\;6f@O
;Ze08B;)S^6aQAb0(de(a.F^,Z^egQ3&H9-,^K<&GX]T\^)[DGDOC^P4)0FXDM+5
?UG0\G>Lc40C81eK9bQ4[3a@a>YU9bOW:3U_)^TQP8-9e7B7UH7U1abCK<MOQgV:
#EU.#@d3cFaE>SUe:?Adb/?c+c4\4+M:STOXLg@cW+O/GC4C/S-X1a-X0Qf9d@W/
&Z5F3aGAK[@M@P>NGKW:D>P@c&V_TQ.A;+4=M^QN6V_5cBe4[7gMg<S5SKg83,C1
^]CMX>OI_f-?e@G67d=M,0BNaN&5)>J71M\fPNW<UJbQa2LA:aO^<dJ:/W87UG^7
dJE9a>:UK\O\TIeCS-aKEO06Mgd3=33S3G,M1N+1#1?Xf2D:DD]<#MZ6L#92cK<R
&3gEGJ8a4#:3JNR+FNMLRO;C8D#YBK&X_HFGf?JNLbDca4WgV8PcU0?I;[+0FVGY
^#_E(.+KD[6XfDO31+IBQ?C87ZfC-#7F(6@A9SY:)b570?)P;6Zcdb18,1JA@g5J
T=#JDaD+JG)DS76/;;F,SKe5SI0;5^ecX?H(=Z1S;UY6B28X;)=<XUX;/B1JYHY&
#Z9\//Ha6BHV+G27-<O;B]LH439e)LB4^BSfW?aH\fa/]+Qc4=,PeY98R.D20#C\
(E.&MeG4&Nd3=E__7=E8>]K(D02]&P3F4VT-Z34cae4]+#EI]54PNa40b(?NNZ?Y
,AK-0BKX1^/4TL(Ec70^c4@2/8QQ5_\ECV\D5E(FK0)RP.>)Z6E(?[RaR5;1^O6B
;25JA)(Ge4-f0Xd<(<5+V-O1WNFe7,JXR41BQb:cLd-BN(9VMgX:c<726,QgADR.
H18-<K9b05YV+S(30P7A&1F0TX=<b&,JH90E1(]SNCF0CZ#Q@Xf4OUDbUATN?]RD
<b@#_QI/T7>b<4Z\LVb?ga+@Pd,V@/:S<^>]FaHd#HRY&B,JSS]5af<=@]8dO>35
O@^Z6^J<d.Y+H=:6/+<cgRB&cQ;<)&5-3^:S)LX-<E=Q?5W99M9D_b5B:#/N^223
=Y_U3Q;If(4ERZ@::Le;06>31AX/]M^PZ6<,;2,9e.8VTWF#/MY1L&4,-TY-#Jd8
]^FF;93GA3#MJb[1G0VDSfLYa59Z&M86S=\VGGG59@?0ZGZM;U)7eL34?0b/1B:0
YEKXGcG?1dd>P)TK<KM6K_QX_M=FK?#R1EM7TL)@(dObX)RA4F(f:;/Fa3e6=]8S
G7._FXC3[T?]e_AP>JM4VEIKHXZB&:RL:+f\:/Q2QY0+eWG(&8\VPd?Z[/6D.:Q(
Y96^g?\-\/0_aS:WFCd:Y?R6H^_B6g)<U^O&YXW@9cUBKV:A<O]VXA\;4,E)FDNP
Web\f,79D#U,e,d0>4A723+/ICQ?Y(MQZdc\4VM0,aTX#(.PL5_3)MLCbTU5e(#]
XL\M=J<a.<90JG_:2bKVK10S9C-4Dc.<\IXIS/0,T<ME/LI<\\2eWTSL6&79L0bJ
CNWV-6)@d\bBTe0(TZIS+8##@.0=B?G<X=_T:BEB5EVLX_=[TeU^G0Wb:B&9YB.f
-Ydc=V1bB\>^#4O>V1M:>b-=B0_,S>_b9N(_N.C^K0=0R0fB61<E],UQW^Ue(\RJ
#bMLWK-4b1K]U6-5A0QDYP5ZF]4:)HPQHAM12fg(E_@ZQR>5d=^/@fLZ@Re:g<VR
=32R^327UGcG19DU;<&O=UV&?J]Sa=-53?5KKcZ?]-ZS,LWP:KLP#5>f]e:<MdcF
&?dBGF1O_03aHdaS;Ua(^;:OO_/K4OX+?6]D:_E287:/?8Z&\H80J6:^;WR@Ng^H
?EdN<3,g91;HV8^9CN3@ZR04DQ.Ha_-ZX=5HP=^@ZB<1M73P3UfBbDXE<KB\#Ie,
CTc<9YZTJ\-)Z0LC:b)d=IgcCK99eV;\74e0TGT7g)Lgdf4FB=2OEWS@NMCR.M-@
:6La.SgL,.La&5f,fUeQY)\RGZYQRS/.F-1Y#QUV;N_DeRPc.X5C>1OeM#\\6Aaa
0A:1HQ;JAW@7fe05)J__=S\1Y2Ge_,CPQUeO2QA.NM]8:0@.e[L]NPQ+TM6LKb3/
DOM6)5Y7JH2gEV]]0Z&29G2?#1cJ(fPda?:3Z7V4]d7Q=c7TcTeT6Y9DT@8[8=a[
F50NX[/@NLR=baAfMUR0J=]BMe;WIF8DgQP4PfF&cV3;&7OO;&T)WGV/1fZM]QPW
CM=(-WS/IL>.:E)-Z2^3W.9dZGdeJW0X=^IEK<C2&J&PH0>5[5N+S-F6fV-F:N6_
?[65<&L#V&MCOCJWO-^S=&^4NO+GF4Yb5b=J.Z4cT<eNA(Td<&B7]@Y(+1/A?FL9
>0W)JSZ/4NBKEg+:B0SY.g^2@eS)XW,=RWZ@0/GERMdO/^HNa;.W<I^e06]3R^/F
<W2=JM76]S6#0Z[gU=[W^AG6f<5>f3+BR\7Tc0)eaMR/:N-06@Z(R5#^6P1(.V[.
A^bCFHdTW2#)Z-[#=2NbDHC#WZ?;G)fOeG3aJ.[&::cIN^CA?Q?J#7_HMXL-?+=a
PO,-HD?7R7;f71HX;J5Wd.ECcTJ8IfK36X]GeX\@=(M:W78IE&?0F/)<0;=QNY7A
GBF@4P@/<.(Cf:.O)R+XGWRIH^/\:QVfa4H058,-@JcUZJHZU@C;&+Y00)\]4K\O
P?1M(Af+Qb2&9V@IadNJ6-Y[&JdEJCZ3UVeXLaRV3K]JQ9X-1)52+.RcG+g@G<7R
^X_#adPI/[M.J(HBK;Fd6\N,.)TOPN_K?/1O+UdN[_@G-N\RRa]/>@0R,U2D^Sf)
[gKE8J(C;XH],59NNN,S(O]9SNL/O<)fgDJ&#(Z.W;@.#WeGdd/JTeXM#Wab&[#;
5V42N^22O(AAAYYYBZe,-[)F=[OFe5DJA^1V6E(B7@K?:RWb=c;L7SL/L5G-bCXe
(2[KD,1f:I(U4Z/a\X&M])-,W.dO:^>Vc)0L1BEXD)0c\JY):=?0CfQN^@;:I^KG
:-cUDK_SH@B9;+Ha_M4I3^K<J8G0e,&O[9.WFZd)J@]6A)7L3N0V87=b@R@TU6,T
YW2Gb;XM0>e;3-&^VC]3,>T.0KOO_[M]:03E7#2ROJ=KVA0HD0#I,Z;<Db3U+Q=6
aObP0dLM?F<[7Q>D7&B??Q+<44WI=\@98XU8eOG(DWYU9AUHP,#-T_bW.Ne30-b<
G@[)U5>d[WHaS>3(RKN^,gE.>/G4f651c&N8FO&f8;&JCU+(^aTYIWg,EPPM(89>
>@Q/7/K0MS6\5\3)MCP_KFIV[e(O213)#^SESB9#Y)LG12d\DYUB&D0TK7^4Q+<^
:5?5TCG)NB99f;A[4F@[?PBbc3c#O.H9gJU]E@1<UJYZ88;T#L99fJ<G@NU._-[0
,@1+b2,&BN<.AVA-VC#595I^=W8<02:=<YRN[<M&d5SG7_B_D4?0OH6@H9DF<eQ+
CHS4?W;L^A-.f7#@MGT7T++MEGBb^SH<]S&4]13GM+.7QH8B<XD0e_>I>(1eW)LZ
O&6V5/UF&DTB7IbT:4EbB3aMIO8<P;<@#@aKNY2JM?_TV=P=dKgQXE<(aH;95D.G
Q>VL0/A3:/H?DW>,CK5B(386/?(.aY(FM)f^CARW]L.^K7/Lg:;L]]7Y1ZEGeG-O
1K]gLe)]Z@D6dKc[5g_VJ&^UNANFNOe3G@W/6Q@Ya,<F6.=gUbIdD0eDe9SP?cDT
DR)cK4DO2O.GJeLKL.Y8If,DMAX#:dOCeDQ2@FAb0?b.R;PDJX1P.CVZdK96dH5[
<&AMBE8OIY8,5W]@8U4E98G1#YB5?)-3Q@R<We.H]QZ\6F>\)R]e.d\g&VHYQ_2)
P5H6UeT+gPPb#I55-,FGR9PT\-=Xg2aEL[bJZTcITWC#9Q=fVFXI&3N9_:;3KP-P
BI8/C(\\(g[G;9PDVAA\MJG^D(^8A<XGHDcfH)f7#<V1Te3RDE,VYRaP#@2,cM7A
A)L0Z+1Y9AgQO:BVJKS]7Z^KK;\_P<21>cGTA6@7d;G@&ea=4#V/.+5>dY9;)C4K
Gb.B;7PO,Vd+CT3@Y4V[JCDC__(FGJY7JN0D?=(#VKO^<82PKS,/c)/F7_O+)Q:Z
GF_P76S,+f)L&fdR:2(VGR[JL)O<Q;V1U=3_[af,)gWf0]Z(2BMQAbW>e_N67U0Y
])0YSSUG^a=/^9T&([8Q[9;Ie:DYK),aB4](SCZC17b>/JaZ_#HRHbf7TEe\N1S#
P<Hf5F0RB>\[LE#)Z):,?6GO(>:<2WZ+1L@E,NL/Y2^aAVJNQG5f@KM>gQF&KgBY
@-NO::.D-7dMOT87KZRMO&a6QNJJb].#C>_,D?^+6(;-bMC<\:C^:g1NLS7G),bH
\0>Tge##c[FI/ZWFDH\B>cZVRdJ)dKRL57g5B),U[IZ_eP0,,<@IgF1K1f-31:NQ
-]/5fXY=/AJRY,<G8=+f#0Y6gJ:.T9[S[@&4S6?aW/_DO8-GXgP:UL7H^>VFWMFP
g810RO#c(3>\0Yc(.;Hf3W+cdg:AV7,FPF#-P/W;=W+fW4A&a&d3e9@\NRI7)L3a
E=-EF6LCA_9_F#B7;0cMDQVaP0A45=;Zb2NAGbV]0NJ&SAM\&N[2V:O)41@8_cUV
UNR0bGNL<)Q&_GaTR<9L:\3+_AXVN-AXgAC;C#f^3M],C[M[]f<;3cI.XM&QK;K+
A).PA)I(5LQW03N_1M@J5_\Sf,&LRbL7B-R,BaEYXdX;TP>#>F;fX8B1L^3@C\Fd
)50=7+O-_g;HPG3EXUU]1&=7V:FTc[C/(@SD+T9^TY&LS^Kb5NW)+:NL5<Pg,^JJ
d]_4d\d:[8FTTeA2+979ec)W\)O@T7Yf6<=W5/N/_&Vb.ZV._JDa.XV8JB>a^UJ;
&eC_@F1S1]T)/MXR3DP\#3HHYGb()eOV6K^\+@-=4;6C_</TYPO6PbaB72O0.XG(
PF/&c2-&d\RB7g4HZ=_KOXS3UO@V,bED[>>&Q.aSb])3=6B6T>,;0E@;aR+A3:fR
S_9,-GQK)LG?:[3Q#a\ef&\P_/,GUIP]N2N.dK73C]/K\8.1KI?)\(<W-&UfAA>I
C:aGP3W8R96C0UY>]8X0a=-170)bD/3LK#.,PFKRAH85_(51;9>g3@]D0<fG;)=V
0C\79#-(9OT7gBb3AJbS5G\,aCU5U77#g:(HZ8WUeFP>KQ9/&H:1Z/;E_cHg:,DB
+@HeL>aUFBNE-?#\G)cX6@5KU3U3BGF<_7&50N8N0_1K_I]D&0\\0\@+L.3BEb@+
JdK#G32<=&^g[/>_g8d)bPSd4H4FOce\[DAHLH-EEF+H-S?,/E-\/&YNEZC8K0IN
TA01PTSURK?gUT\1=IXV))6Z4M=+AA&7T=8=_=W(#\;696E5><@5aV8Jda&P((d1
PPZg:5+36DLO7-[6<1=Y,c.QP^M7R(/#R3EF]\@ZG68SQ1DY]HVJ-MKcF]:L]#1R
gA_eY),I-Z9fddd6K(H-[:5UO4a.;>_P&9aK5)Gc(+L\D:KAP+(Xa=<bf)Td)fg/
<&T2PA&-Ud:QPM#,;FS&^N(7-?2,KSD?K4R^##P;,4\Ha1^DKCZMeY]>R=R3bXF+
O443H=,2e(W\#R&^=TF#GKUHB>:Sd><&2(KG7/dNLOaSCaLA]_T-F?R1X49@1Z?P
Xb-ZR-HMA0)8J8N/5>YE\PPYTLU?N4BKPGcb0MV1?W777XXF<G1RZ&>aMY7<(([S
6V(XMB)ISa<YfI7[TT#e6-+#_3L,)8^MU&\5Df4K(df#L[Hdg/)KYU-ZD;AZX1Bd
YQ]9H(AQ@d^ffdRWW;LG0-TU61Pe9)KZ2(BH,=@M+J1]RfS[RbW]ZB88+e:;I:K]
B=^ET]9654J:?WTLIB81X]b0/Q76.d(E+]H2677:BS[-#72&4D^L<,I&W6<\f@CW
\3A>Cb1N#Jb1TGEHD?7Z/^8XJ.\,]g(PG0.[T<eC55Q8J8KTBJ.=]-FPa0;R,#O1
Ta+1e@)6[>+C0/GMM.#[8R[1>QTXB)f]\Ug1)P<O@+Q_-9I)W4VZHJIcZM/aFI9)
XBLL9e^PBH7@+6&Oa#R[]76B?XKPR:C>P-^B^)G[3#a-N90[?gZ@I(=-85>I3017
_O\+1=727,(D4)N_+_Z_;#R5>+_Y)+E+#,R\>O1RT=YCa_+F;KBRFI2/GL\YX;Ob
W@9I1R18#U?QVV3A1-G-^Xg_W>#DL.3A)M3V]aJ[P+(c1aN+-9YNZI]FG3@#OC;Z
@T,[D3Z7DFW<CLDaL[e\_G-9]aeEJZI<=[.]fcc_]eKKAPN@_Gg5b<Q._2;]C+CR
?K4#Q29IZ(L\Ig&-aT#Iae8A);eeRIf\4dV1UY,d@>QeU8KbPS5d+?PGEe/aSgae
X71^73^1RX9<B@1d<(D8a\?Q],TPBA^S2MR>^UPgKUB<>BJ1I^96g-9Y)>=D]#S0
RUg?-\-V;WOL6HE-H&_<,WCMTbf(7]?=Q1+XEOa#MED.H(N;3RbDFJ(M\L-39IK1
S;>J3=;XMceFgUdcL2LggT0S35@+M9SXaY43NM&fe7Z?Xb_BY41CS6#ZR28.KFS;
+a(#4F^,SC5.5M]@O8M31[/=AEK&TR-1K?Gc,JOEXW+d=YSKVWaE2=XKR=dW=,^/
]EGM&JaE\AQ?L[(XZ:,J(]H6=G2U)=5V@@Z+#9117F\0:#-d:f;=?a\f#dXETd#H
.D^8?d(7BY8:+eD.A(/S&(XS(dA4Z)L:B+];e-+A.J1NeH@6:9<8)PUQ)9GKU+b_
=R>]#;C?7#V;^#AM)A^X7_QcSe-UP^)\A^.BgT,)aB<V06B6I-_:6WDCK_Rbe@[\
>HR>b]/A,e+c0\V@2-G=))8\879P;BGe?-/&=H40[LURc]+8:XcUT5DH14YS&X53
N;/+TfL6NJcF[U,ZJ7,QfNP.\69dB7_bc(AO&7Vfc47E@:bK<1^,:Z>>Lb0@PM6C
A3>5a,<aOf?-(e=e\e5-H@#K][O6/IdUYAKbZ3Ga=I,\RG4g1H4.P8O@;<+;:>.(
8KV&1(cJZQ36[ge,4W<:MRc-XKQ4#H@[>+,DW#FH^ZP?1I0C3#.,OHKBI)3FA_UE
6Q<::JI<.0YYFR)4L[OV+GZPeYgQ^GXf/H7e/F,BL_D1INV2a)O&=:ZYdD>?4WVF
8a2>-25WGKJP2RPQ#4(Q=0_b#1,XY6F:,OVeHMZGB57-/?D7OG1ZIaLEe#0;Wf[:
^0YI_/EY[A;DSQZX.-UYGFX_NB&J_de,R3:22#^:.B8-IbS/I7R9L3V/;:H40[b-
eVfP&=8)@KB->=K@PVHO2ETB3^ICR/PT40e6D;,9DQXQ>:8/c41a5Y4/00Fd_8]F
QX>JgB^R>45RK80#-ZdeO^?BbAAT@=]XB(0#5HS6D]].S#MH6]B00N^+/Z,XK>W8
=YAZ07,^>a05Pd78013=fZ/.J_@4ab8KG@#H4fLaZe06]NP2-EJ_5\3U/40#ODKI
+dMdR[C&?R85dg/H[XHT?8MaBKCFfFVA>d&7N+XR431CA#)T<e0N9&f9O__dBM<5
VL,_-BK0<5fE;T7,HE>.AECdb6\c^J,9).SbE^-MP8bH0J1?2@;D,-Sf1F>1X>+^
8^BO2#LP\fDY);c#=SAXf_AW7JB4E23d-cgYOMe2R:a]Z:89cVM(TW&DEORCS<K/
?]CaMYNN?1M55fNX-aIgIBRc9e0HT3/VdO:1^T^AJYb>,10.NI_YKb_LBfZNGdQI
\JQ0W(Hf+7&b]UXB&/;#U?R@P5c>=\LD-O&M2TXSHN@2a:C0fb(U;cUJGa::V7:^
dP+#0X]/?N@@cd/5W,-\MN8+g7_8FNS+Fa4IFNO&5M[?3JOWY<(g:#?QaD=TTUf7
Vb@/P^SA8V<LSR05O#d:E5)=d4<J(4a&AB9b7I4C\.b0NK[1]R=R(ZJ<1C5&6=L\
:/,YGce.ZO.<G.\EE-?NYHD:DSI@dMK2+WOCDeEN/U45:+a;N&HM7CKC[gLR9+P;
\NK=Q8b\ZcB151<CDgT-XH2>Y+&W[5/D6[UW4>3F6I0MJ]G8H,bS8]VV4YV+Sf6a
:7WAC]ZT/+:([]3D\)DG36cKRW]dg+0<+]LX8fPM@>WJFWf4[B8K_>[-X.1U9X9;
+gS?UPV^[Qg+\;U3?fJB-a&_HKI+K]]NLeAcbH)?VLDd/PN]AE^)_g:^5K1b,bHO
3@XFYTV4<L+]AF^/MT@\c<A.Y9KXEVA>1G4S+M.a;OP-dSN-Fg=OLZ]<]cU\1S0Y
<LA6A(eee.59=_ODDFgZ,)+[DGJ;e902Zg=[f\e_g>(=0\>4Ub^+0ZLfKVM03P,=
CDAd87_\[@Z@bN7TP]ffETR-)[X-9I9;G:?_T4KdI++EPg6)-4O>3WQIX3P272:W
e8<L6DTP7EN40M@W&@GB8=C:96.&5c<<RZ-gP]8J-=EDa[G#Q/Abf7gT?5&[dH<M
G/]f+e^+f)AINZ1J<S.E;VM1X.N&;Z[T59Ld+aGR@0L-/ASddX-][L#5Cc?UH_^g
--JUAH5X1@_R3928F-L\gE>^TaZI<HNS@^Z6<+g<QR)6=61ORD4/L0Y4BUGQB=NU
P5\X@\#5Gbc+@^T@4>=J1TTG4AAWF#+[bbFD3fK<ZCU73Rdb?eX[930^)cbQ]JbV
@^WU>gQ3D/5+IH1>Eg8+d3cR8a?/:aYTK7\[4bY-O+4.&SMVB5f#=LXK/_^4;62@
&d>6U)G39-:Z[P_7.13CRUDdXYOBJCN(7.=A#/dIF./89CfF?G\Ng#0+&KZ9JT^J
Rc2C8@46#L\&)R#4Y37D/2<DX;F@;#&+dQ:\_UL@HT:D5:Q\c.9WLWT2Hf?aTHK<
AZCLZ7dT3QA(GRL>eEA[#>M-d9CN.2#cE>MFAa+NG^Y,[]V6A>I#(R^N]@UATSee
U]G:7fOf<]4XN&B4QD1D^7g8SdRUIJ(5J00LM+H]C[2/U^>0C,SFD2:Y5>[H&[/Q
,B>g19>XV[&c+DGN1[^K^4E(]NJN2c2cZ;RGQLDW/C^7[NN16L;]+:2Nggg\2V/;
RZ.>J[WD#,gfZH\_dM[J>J&bUPW/)_3FMP:f@\C@7\0\-B2)RU@CZCHYETc+60)X
9S5DXI+WW<g\=ZJ=;S7<\C(_\+6d,2(^N;6+-L/09I;E(9;V#[ZU6724\;ed=R9U
\2F[<[NZ@TDd7)_S.\LK[aQ+;U;,YW-U\I,g)L&E(5[]g2BTWcHT^OZP^5K#@);6
e;.IZeb,;_43:JU(aF_W4[IH?&<PU&N(R6&-,YAW,c6J3J1A\]Mc,f_<#-,?KS&a
4\_aW/&<ZfN</[a./IR+?H,]+#D[UOJ>Y&e>EKV]QEbHK^^>J-)dJH8+D+@SM.<5
?AFGcbPS6a4NCEA>)/LL8ge-LI<e74N>OH//J(AEaV?g^6aYRFEWdbgO3QJ.-K@W
CWbd3](P)JgF&WB:EYQff-VMOWJZVXCOG/Ff+2IeYJR9@_4dgNZVH\Zc;C>V<Y_?
@UY)P13LY,4(=)e6L<NVKBa3R/-gG&cfV:H+BW#?X>f=WY)T/d\]_RY\VJ#4)S=@
;QV#]ZK:J]GHF5W^:fTH>?)<;ILa0L8D<#Y\;)HGZ+-.W75>?4KR/UDb#:b>FU+)
Q43@9d(T2Y,<#@EH0/Z-E7cI4cSa8\eIF.\+6Y[(?B-\VH16L@9DHQ[.ZY63g-/>
P,B<Y^(YO9]82<1d6XS)I;#f(:;#.\gNETE@b1g[AcPT;#gV4d&YE#a3[YOBQPe^
KT;X7KSA8?Pa<eL<MbXGf:B/+\50VOZ8.I=HDJ;^4ZY..B,ccX@W/PV([a@U^gZW
>a5UTU(\T,T[MKC4DcR;/AW4BgV\[J_<Q>1f6+SIU2TKffL#>.VZ[\DGe>cSW([@
MT3_:#aAR[VIQKbcf/I>7(ZeH8#NCdOJ>#OP++M2)HcRDf]Ug?907bA6J_c[^\F+
SF->044LK1>J0<1O(&b1T/ES,TTH]VMU\1WE&#LaT9NKT3]cDNg+e_#O&[]9gXOf
#Rc/_NJULAH]f?ZSWeIL9W5_fa@#-[(./4]^V>H3RBdQ(R>Y/QOb1JU0S#eL6IG5
YYRE\#,7ALZMC]KbE^ILC?80.8c0CR_C(JU.PGNG/;X1L4GCPITg^=5<F0?E_d#P
N6J)7(Rf0a9>2&BYIUBI-PG]T4.[48M;EMdYScKKSdcUKL7_[MJIB?AMU8/@WP-#
I)MS(3YD1F1X;A+Y@YL>0R@X3A7Oed;]X3[=@#5;5FU+SLa037F[P6.O-^8/2ANf
9#4J1bJ+Gc:^a/C(CQZ)0^(_9V&_\+_VR]]#_<-]3?e]2ADY];,.F68(AXGLc4eH
bIBNK4W1]_AWSJ04/W/+EZN7:B;_ULX;+)DKP+CB895^R<e/,I\UG-e>_a;EM=W_
KI7G_/0\T/1K)_a@8RIY\:\T[^aF_HS6IDLLe?g4RV5QFF]dgK[+g@8Z;IfTc/\_
NF49.,I7RcQF3d:48>cKO/0E-9eI.RK0O2b]b75LOZ#\U;,If/\-RR@_J&Q8Q210
-II((>A;S0_+;TN0[R(eFD3U0@?bF;<e_V>O>=Z2_D@LbUIg6WXWK]VBIbCD;SE=
MGVCXFAfKFO9R:/\(IIa=Y1VN]7D)0d_TVaL:MMfX97bO/=O:9;ecf;WLQC7C.\A
>eW44-7f;a<Z&L(JLHWb4Z7WV#[6c<OLI\=U@F[U@=Od=93_=:d7>DHA9]/(T=5K
\,.\SU^>d]aV^VD]=5Vd@3->Yc3.PIFR>N<+PK1da&KKUR7TG]IXDPZ\4=M))CDB
<F@RM9D>fB/IY1BeX[M5O,F./06+8c)Yd2RB>W,SBb3^=_b7S(;\8,d)12eIL/,^
JX4P-6Yf480\1^0?(;KV:4D5JCf4]gD759KZ>2JKB+GT#MeL8:\CM&eGB/Df-UVH
5-;P;f@U\JR53Mf1\3R[#Xe[EdR[_-<d?T^_O^-TL-=.3^7f++.a;b98;,FY\a>S
8UD&Y/94c/8+a@\.\5L_Kd:bELe#X]@DO4_#>.,U6edA5.JJ<]aP@<SF16GWa7:4
P._BgGd,C]>V_=LAJ^>d6<(6e7/6gCcDaZAFL(HQHDOQ:QR.)-C3KKDWDaR1C^Z[
_3:^>+4Z8@B[H-QO0)R1e[GCY?N./3_@<4:]+NBH1[PH41#0+OYaMX37@P[,.3GQ
T?R\;0&74\-L8,>G^^K:R=_/W(5C1[QZ)D^CW7NeFgSRVHV#=dbN@?EB8VaY\Z@W
E)LC8S.B+(HEZ0WUcb(+^+?BWY:E:S/]?FPCU#;(aFFAG3JJP25eC=0@L:RCg14_
O52@L.R,:.N#/;Ic=K437NZ&bDZ>].=[(VG,)?ZggH[b.4JZ]@acU1(K7Sa^S3Y<
0Cf17M9bG6L)_?G<RZ8.D8Cg0]Z>^)D<6L8Q4MAKHeHSP.aBCXI95W^9gIb.=^;2
TG8V@^F5M/b1T?.>a>Lg7L?@f1^HR>O#&QK7/3^c+6GAM@:\G(T4JaT@8V[EYV;_
dLc/^Ge7SR>.L(g_X6[_Y^)/7RV6Bg:/IRDKYJ<4_O7ebd(@U&N5I+g]J<FXQV.)
[,A3OMHK0N;R.R8&-T==W<8T,ed5b),&@)ff3]RB_?f9;;JPT24fGfH@FC,-U8G3
(HZLH8B=OVI9dN:AAMEF/K3S-Fc&\[+[Og@[^B++(M6JFW;=+BPM/62GgWDZb,,R
<;O_P&bIJT\8;=]+PgB?=AYEMRM^NF_2<K?P+U2]LY;?S_63@gP<&+OV0XKW/P4\
[CS@\Le;d;7@55Q02F<(9H@7F95IJ;Mc@SbRLLZ3K0<CdFD0TDIJ<?(-6F79&KTI
Y=0YaOSa]D?AJB/)PFTJc^[E,XC)9KS75eT2aGH=L^RT<aQ.=AcXDAg0cX)72/Ye
5F0_9LgMMQHMcS=\;dG&f(&.OVKLK6E?M/BZAQ+0^^>2gD<V&GFFd1fYG:M).2aY
gKD(+\+dL[JDFD[146JNJ&NIQO+LE\GE-ZgVKI7H2-a=;94:P5]F9OAADM:,2.>-
-W^O]<#=9?:9S(MY?]eZF+M0MZe9[K?SHbR[1>(YH,X>dF],OQ/=V>F_1@J,?>:4
6T7[]LSSHJ3F0L8V&0Q8IU@N4B_34TZ=c(Z/L(b?4<?=a1UU4F_G:2L;DWP2=WQ7
=3Z3EY?SfZa076YOLTO;\.&BWL[^F7HV/^#5ADbeeOa[]]b9&7V3V-2M&B>:8J+Y
UA[FFMFT/FFY5GP^(C0F]Z7Uc<O>JOIHH3Maf7QdG2O/\g4DZR,SW4)HDO,L_@GY
U<F5REK:e[=A3+<.JPcB+2+AIY0IQE?d-J02&QeDAU9,&E:=GIAE\B:aR##KLg32
WdWGKfDITc/YAOVN4IL.4:S[0bHVB7?B8)7C;a0-R)bG6GSU1RS(.8_>UMGD.\KQ
L23LcRWE\\?7I<2(3geX>+00CPA.__(g:OSPTL;CU\a=47Z&81S\T67NZ@:&_g]g
@Z3a[^&#bU(fHCX/J;(/BUKLPUY#g?Q&Va1/5LR>]cW@d8O.H9WH(KH@.ARJU16U
U?,@QWS6WF_f8P7U,H^LUESBKV[NT@PaZEH9\DZc+(Y9&[UJJ9T^GQ#:BS/#G=F7
#8MY3T[5P;+b5;)NN_E\>D5_\Vc0@_LW-]<W=QG9HYIF(VVX=>^/DQ,C#]=@4:I?
)Y6<L]J8F96?,>VQ;F)&HaY?:]V..^eFJ3,a4cCe(6JRJQZ3KW2+Nd.H/,>->87>
;Q,1fCf=.Wee<WbBR)=2=@0YV856N>#;#FR)J&eF;3f(=.S-A_2CU)VE]@0]A-R4
R,<Q0PFI5J.\&=X/=\:=g1GJ6#?a?AT@,[.R8dHfLE+O55F2LN,^-NLDA/fBH@UA
gIL9C3_E@W1M&+0?2@./SY50#++8LI4SSPS,(YGg)Rc<J-\/?>IFK6/J[J#8O/M4
3g?US+.<6/8[U-8J)-<A6M2NMVV\XdZG0g1@+@>Ca(VeE]MX^LdSb<TLbI8/WHG6
D\VJ).\-G-7#?Z>9I-YWW+3R@S[X@LLXT5L8CL?M/1FM+ONbgDHKM6I(O[P-V<CX
N(YWdfOd_&G,&64?^HU_HW9dD]Q&S2]N@6@\J(;NKN^)(..IXAH;F/W,2<SbaFf@
Dgf2?T-WcMR5WBBfUP+,b1d^G^e)JTc6O8,G,TU]9eSS5Vg4/O?Hg-<K<83<,\WC
./+N/Eb+/3>/20<B]2_LCaAOC+8K;6=C(Y3ZT/.MFE8,J:LcCcA)d,V2?T:4-6Hd
cBPbN^1d<ND9.-B_=2.O6fH)=_Q[;c[88GVN+__QBKJ>X[e>Z\09V\KE&\;^OXL&
+Oa<K+5>gCf4Q18S4@A]4115?dQ]N[4X,(@eGg:]TSa]bY58/&:-\Je:SeSA2f[G
RP-<gEI3.E<2XEJ[&;\;-433=Kgg@GZJ\W=?b,-:I?(Gc,:g\PN?EbQ1,=+d=#VP
P1OMc].7ab4e2/Gc(U9V\04Q7D?+[IQ36,2ZXO]F/Z@M47gW,FbK11M,<5@U&6IF
#A60FbE;81B)Z/c>T-??&:)6Y/54)HQNMd5T&I#-D(X@AM9=3P\W?\]0.d<e]OFJ
(MX0HNd^ESC;Q,[;DF=&\I.@B<N]T;QA_U1;<LMQ#4.JF;.J_9\)+UK[d&dJVQ.\
gW7P=@G7(=DdV(d2F&E57a6J=MI5V8CV6ddG6f@)3DL4UE;Sd;8egAdHOOVHFG8#
BJ#.&U;#(^>JbCE)+f[K#1^B[6DB8_(LY96d[10fCfgd?dU\ff<1X;7MLA^5H_-9
LF4.Q:Z>WUg4V>):)6L5SEMP6J8=M:FN3I_LO=ZX-4_#fQaFQW[^&E\FK)S&?11O
MHY^=TW,S0E^CL?\Z6Id2)>-.N=NdJdH2]aVa9<b=RV2M<[Qg]0]=[3-ga.VCAUG
O_=If:C=Q^e)&:5+DL=&)e\[YZ).fXa(&Xa:VDKGV=C9Rg1Q0M;V:)SZ^VI<e/52
+g]NX=Wb1/GU/<30>6=7-P-J+9X]HFB?1<Fd3L)VO17B(.9EG,JRI?>YTDg/BRJ(
_C]9=4JGg4aJ/ZB@BPN5@&LFJ^NH,IMW/bd#?5QZa^NgeCWX1cM=U8&O/Hca).Yg
#@F7+\=F^ag0BcNYS,-1L188IWB?g@9@I4=M6QSWMCKZd[>#U7X9#:BF8H1HCV8D
YTT5=3V(e\?8_JE+ZJRSY6G_3W27OY@+4#E)#SPVDSd.<WJMKfgT,eXHK/bF6IFB
55Z>7Bd>7DZ?O(e0:Cb)_DR;)]<EHe)?Wb(F5GS5WS&X54^adE-LJXJ+_9d572R=
SKA[)=dKVMdHUN>[GIGQCeELW20S14R^FW;XN+)Q,L:Dc1P7UPI7_9GNea3HK:F-
GY,](O6:\,7b7;B8+MMH?R;ffS,->^)0MeEQ,QF>=9Y-@9U#9J;5W-.>DJ?X_-#O
>@84(BV;a;K_fI6K8V\/aE,9gU::LdU=&GR+^Nf(fQIc/>d#DV-]YGG8\UKN2T6;
VBVb-9._3TCG4T&DFQ+R7_&8#ETXH+:SQPG#<J9LTRYZOGW8=#4JS#0Mgf\:=C4b
)cK>+dN>fEZe,4N;K@T0;I?.@MR_61>:^UKgg<4.VAd?7H]PPML(/9P^,S6T8CM=
E2IA3:fg=XEWE7IGf+Ke=9,^_Z0RSV=J<QCSBCagPRa/:0V6V1PcS45c&G8_g5OZ
#1&Q\PE3Ggc]aB6-^?)/dL.LcdI+^@XH-fCK/^?\5,JI==Qc)_8<Sa.OUW74M^Sa
>eOd#Ug74e4ZL6,@0Z9AcaJ.TgRLINQ](-E,W3_@aIG(VDJLSQH7N)&^=&F#G^.C
OJ;>&H^UYb\WCgcX#.XVadN?:1_f68e7)f[M(V[-5&JH_<M>R03#@;X(&3XNNaJL
-+N>,0;YXBBYSOdJ(O@^A<@C,Q+94]6e3BYMCJ/S)J2-\^=9030Qa;eG;GB\BN_,
6bHaOK0T1H\5f>^NDe<W^HV;6QOa.)dBE@Ae?4bd^T.C=7A[Z;C]5K193?eb,W:R
aaZ8FdJ/OU7OaF.dN8M..NVW<)_0-ebaI+=>8=?./1Z(-JI<FbWDCgRbJ(,BH,ad
(2=)M31US&#<)9XBJ@A/];Z@[NBU;?[LLB381g;7@VHSS,8ERM=aJU]>(<UK1N@a
4/>S\&a,CLDB+RAUM@JVfV#D/\=.>@7#Qb@IJN]X:e73-<f)#V9c57VNE2W/UN?[
^4a?2+]cHJ5Fc:V9I<,Z#HPYANY;)##DUR=Q&8+AH5Z,X@LL4fW<5L;TQZ7[<P##
4E(T.9F&K3b;+.<TS-^d2XE:<aMS_/RIZ/Ug;RgV3BFXU)bZ33a@fW0gUJF8@H\C
HKM(^>HQ8V+GK.X<d3G(U9<7Q\4^_\fbLBNRBX@eHg_=Q_,f#;b@bbHN=#AS1)eZ
/V[--Q;/O1BLF=OJ&NVZ.+eF,J,7Q7+<CGW8&L;+04<OYg#NNNHS4U858;<4IOdQ
cO+G]KLN(;8(X>PHKMRZd@@SS[G7Q_CX0F:J276\:ga3_6MI4a\D4_\Qe@>2X#ZV
J(S^dT3GKdU2GI^I]gg,=;TM^=]3TC<BXU;[B.U+Y6W?7<7,@5ETK-RS)+IH]VA)
4NGLE-8(=3>I_fEeS>=N.eLG3FAP9Q7&-JFBb@R62>LY9]RZS&51A4CW5-<9:J.9
&-#7M+,P-U\2:)VWP3aa39K6DBDS,+R\Cd-92?Z-0)<3X:B4[#Za7O)TT(QL#-9+
JJ<cWe@UgbP4c4\M_EX2E&GUW^[a)ZUG6g7S[EPXTHY5<Y=(P)a?g[Y9>Y\(W?0F
_1Pg#M7Mf<\HdK;.XJCWT.J7&=12e&GU8d,2Mf>1ff(.RS>33AVA.(OWdYG<0WfC
<)TA#]d[Z.J21Yf&2D)H1#fHc1D3G^&3LeEW^,[\4#H9\+\J93?GN[9L@F0;3+[/
32)-\g)M,;KZSfO3N[Od+S#5gP1HA\^YHdP<bLCEV;Y=P4\9#GDbM]]#KOf0Nc,J
5-]QE7.E3beRW?b_.Z>G479L,M.?Q-59K\@gXK;?@F&eC:FDHN-(-T3L_CaW.21]
_3YEb_BIPFK5/6B[;_)3RK<ZDU_PH/+/LZ-GE&L)Vd:6?Hdd>VP4aC>cfbZ^61H)
RQ7[aNfT0=f]G_dCP:Gd6=XCQ<OJ[_H;KBVKV=G?XU3;YU]W1LZ0T#INAdV@bQ(M
(?P1RSf&Q+4B4#W=MVSAT[^4dFa):d=36gQ5:##J<F2FZIZ@.[gXV4=8&DW-)9]?
,PJ8,==\+b<I>0H(S9cb9Z3S]OOX0FWa7(0J=F.d^,gZZNM)?:U6@JPdZe<M4.==
+-\?=:\)aeF(\EZ6K53:g,T1eLNZ>&6=.+DZ_(A4fA[@D5)YG&8-W3fL?dU9f7XD
DHQ+F[.d^TMa6Xg-YggbU.SLU&[6>4N<=G,LO@>G@c7?7+=.=;cEdZF\=1bV/KS-
_U-KAOC3BCc:AVR3QbM1dd<._\9^O]F@:N/cd)-Y;]d10/9SEc57S\Xb1BSV=9BO
I1_16U&TcW^Ag7dU0_M[T8=8]AAbB+<fce4/5eLKXDIS#YZ8fO?cU/dIZ4B>@/Y6
<=BK1:g[Z#K-A6PR7I]GAZH;W^A]LL_\gV]Bg4(VBDDW4&]3N,bGL-@O?W-^fL^f
WZ5WT-:JO[LadM)A2E]#[fX_^?4S/]Af4IH,&097JAIKZM4H]3:\Qd;IJ)K<9#0P
6(?d,b.M>CN0-+H=4S;,&YHF#/TW0H_\He@g3HN\#a0WT/IN/#J>dX6[TA^E#AK^
-(7H9&3O\\[D+;=J&+141HJ39&a?O3]((M:8@)IN9];.IGeL0(F(e>>_2XNecaaE
7@>^Z:6.JJY3<QJL5B;S+cXUH2)g4FXbO(gTWLFGe;//X2g0VPEc=?./#gW.>I90
@FO_Xa:XSG@8WR5b4BO)V/^G]E#gBFT(9b6dZ>4<[>=9^EV/2B(:7eB(/4S#fcBe
8-53IQG7D1(N4>55?6H\&7g]A/&Qc3\GYTBV</XL&)c]Q]95,^:gLgg9Ib(H<JZ?
dG@;I.ED0V,QB?J,?_CWa<W-)^=P><dLU-V-?9D5D7aU:2..0X3(gUG_3<[KLQ03
eU]&WKHCFb/aVN>(^/De(NI7SDS8W#[J._(NI6O?7&?f6^B9L2WA(<O-(AKM6PfL
1R]dbNf7G(Sgf-M,SW&.UbF/014=bFW/#<17D0,bB0ASB.4/Gg9,BY=:+XAT<-8+
=>23JA<.aWZ7<Yg+C5Q#PCRE^e;f4M[4/;-GB=C564,8aTgR#C6Sf;?+VEA-V@P\
2Q:G#LRUUBTDL^=-UN[R]N;-C15,XZHM(KA^Q34E]\^S>EK&5aXWcXfcQ.9V=\8Y
+cS(Y^fS9=0XbB,3Q,DL1\Y_fe[_0:f=HJ(58Yd4Ha+HB_X^#>e,8L6(5>g;P#=(
IfHK:0+#;+0EK)9@6CbVX4=fHLcBX1TEUDQd/U<.E=(b6@>SgcUOO2)#LRVBJg#+
A>Y/K5,-O<B@5T.:M@Ma@+6@8]]4IbR;3S1Q+TQ8IgcE(LNDfWMZ-)43dW+?Sd4;
[/XMNO(-f7:YU#A4NdHH,f5eY\-//@SCLCbZZSJaC8QD(>G+1-=3g]++V\g^\A<J
:E(+e47fdca&/>EdVG0V+U:93,R35@&.DCK&8:U0=C4JG0,@/E>ET0N(gJOQ&74?
J8Z(@=PcT;3)\]W;SMPB@K;^+CFeIe5L3Je:2LB<Uag_H.Q6;=I_3[@+eD;;J6>>
4U\CTf&&Fc(OX/_L:bRBJC@ZSN,_?T>XYACDRI^ZP.3-]->QWKfQOFNOC8EE=UB4
0&Z<Z#XeP?.SO<UCI5W6dJLL&5N.H.\3;,=2KR4\O4B7af<HPY?[G30OC\HgK<OG
J@@4&([?]CaJ(PNCRYZ?:S505R4CZcR4:6DfFM2N2<8#2@5c/ONTW7>[a&af7,U,
NTeT>;,V,?H,[^M\BJJ9AQSd907VcG(Y9\Z;__LN@TaGK4g(4@U[<6U[f<:@Y92W
4b5\/#S[(dX8<@SIX:9MC:8(YQTI()A9S+_g8NB.S8g,ZfZC1_G1a7CB,,^9L\_-
YELX4(K/XQ;=AUBeJ=)c#HI3CPdUCg:KRG>a0KOTN:/X]]&##YfQNY.BdR:QSU^f
ac&]0G?1gK()..+\#S;CV3Y7De3b6VUe61^U>3O<,?WSSV/NK86\#c?DAUV&4_40
Ia_M#,#M8]FIVZ(E6&a?^0F@JH6]I/UYaC)N#gNY[ZaSA<CaT)7_;^ZRZ^e=54(?
WJZ1]Qb?S1F3dF:<F,Oe_,>IPV<72F_R/):UG,R#EVIYL-XbWS5X:5&OTSJKA_@d
6(aJ3;)<S81MD1BV(5KQdAGT?96H^Q=Eb6824J;5<.@)8:>SZBBT1GNJG[4KFO2O
CLMBBb,4Q@PF964aa-P[]<;#;#Sg5T_>U-VD8R-E2c[c@9b8]=[_QLUKT<NCVE.5
_AO#c\>FK6JAgM:2QC<@S\5R-OX4(?ZS[^IAG>KSQV<(d:a/[#_3[TGA\VgHg=Q0
1]a@P&A9a+8.GB@QNQ,=Z?/VEEW#K4f9I&SM/8<4-K_dId4YK9=XW?_g6Fc7:):a
.>]3I]S.H6V6a_0&c0R&D2SCX0g<V0,0F]K2D+(B<L<6-)=8^JT1-;3/JZ;R#TZ+
(d8gK8G:_a(-)VX/8R^10Q<&bENd?)56;Fa\V3YMVDTfg:J_9=9fQ[CUSX5.<ff3
7W0FgK]GK-HMYQ(79@JHd5EL+aEe\ZK2K]Kb3O=6fbJ#P#X)>SK]4L=JD/+CG-gI
J#(+##1BALe]J.0F,V]][>A(P_^/Pc3fRR66e^T->V>N-P]DLc/1OUIT>;?cPFCU
<_)(#EG2T_^4KC1A)^R:EdKJ9+]W:#AI\(KSE\V=OH8(5bJ5:E)186=S#7D.T-IA
Ad/UPIAP[)L^a7]aaHRacRQ^+W3WgSD3Y#(V:LI3.M4NJLLOT;=BYR.MZP:+>MIf
M22K3b8-e2EcS&c+7F/P+8J-N^O[LLVW/.R[3F&J:U#K#UK?/4)CF(6@(-N/(;dW
FTXTRa-3E0A,aOL9NWS(C,F1(UAJ?3[.:b.>YEg\[2,ERO[/U&R::MY1:4+TC]?W
_JPT;[<T(L3UK3gXd]^&45Y1f2;gf_,&/98H[=4c7F9d3cI+E2e=#W8<7B571,.^
-#D07&SOTdD_LJcA^_G)a&ARff[C:bOC(-Bg(cM@gJ9<C\6^ZE7Yc6Y:HH,b?X3,
U=@L3&3Q-4[RYFE0^7WP/47#P^EDIa2E[3bQ=3_&T2#CVRD4HfYdCA66RWC3Q4&J
P8-1>G1J-_=G,RaFFd1E;YV&-IXO6N:M@e,:5Mee.Ab=2_0ZYA>Z+5f_3XU)3SFP
N7:GeY1B^S.W4@,e(NOSIf&WP50(Y4OO6V_N;QKO6+CD(/.;85G9WM=/HKUdY,4b
9_K28D[VOYY0-Ua?.Q_A=>DbIbf+IXga.PPb[?>[,gO)bQS;V8GJ?^JaYV3LK&Q\
S+Ma3dVIePaP-HLPa^,LFb)]7Z]8FSd+9K,<d+XVf8+Od^1W(<TU3W.<-N.)\(?g
A6>\HW6?/TFL;@=V@KR8^3]->/YEYJ)P\S>Ef34T+FAT-:QcDN7PN:)/MTE3AKU[
Wg#0B9S-])^V.1B#C=d&PBa(:c\__KL]+,?^J,;S/],RT)cK=OUPILG\N/Tf=8C2
?D..+aaVPEG/A9W+fFK>^<GBA<8ZF,#::LX]>FXW1g;K#c1=1KUYXd>K5dAM(VB=
U38H;gP(0g_\W(@b]0KJZVORPCD&92FK.N(^A_RVL0gBA5gE3M+S(E2N@ICXCV_<
Rf&2FY96_B?\Y7@[68(Yg@Y.8JDL/H?P]E(Ld2UX(<,:WKXS^ZSS4;HJ>(M9:R-N
>B)V;LWL:[X2A_#,?-QddgN1g\:bTQ@dDF;]DUaR_JY#0Pe=[<+=#8Fb[0F:Sg6#
#Y3c_X8R:Dae<bEa:TWgeJ@_#)#Kgc9QN8B^S)2+OXO,c;COFGYPeaT+WYO2=]T[
1_KL2&WB)f.7^>7\\cf(P#46W_4:,FIcK;L>;PA4e@7JDUXV+^W?WHTAGf/6B,H.
AANPV4baDP0^^AD^1BIX)3T9Q4Qd&PBD;-VDBQDQ3)fJ1BT=CNPG;;)W,/&;&GRW
3g<&_E;ZEf52,RX+AfMbaK/65(X6ZY))<]912:]?]b->Zb@<P_d,1ZI[c\e=Kb1a
R6>[CV/@RGe-TON66KCRd=bBCZ(FM]aG-RA-HHZ?Ff9<fJa4/M;TOMNS_SP^J\)>
2#C_GTN&J6-GFe,L-^ZY4MS,=/@Fe?IG)#:QBF36@IG=2=V,BL)4XF/dJGYFA:#f
8E:?SOG;U.C4F@J1KRS[I_L2OYU8LWbZg#57M:1[2=7-Df4^e514)@:>e:H]+9cU
BZ:HeQSW;Q-d763L>FVK.H\J;3DW/:YKH=/)[=9HGG)\/]U,UJZ[(:DF,3XfL7X\
UN.F,U?,BbEU6=d[/fY.W;0>WN:I.I79\NQ3ZT0fV&;_]3&_e#CW+MD+69J>+6:^
SR1?/T9JLQY88QGV5NTB<]SR7TCVH0?>fIE6^OOLa8OC8&c0I40UC9=1(G2E#(C[
&QT6bC6+g]YDa]JQOOEB-cJ2MN7NXBF:2[:e30&Q6KN(V^=PDXF4,4:ATD<ZIE/G
V):Y#XQ@_P+8EE/OdP8SX66(-&JEPU9E#AH7=\:ZFgR4_FfWXA3YRH=?bRC_QRMR
a0b,SEGZbd/KSK1Qe?S7@YV;GaMOJe1IgL2G>gG4b[EP3I,M&D\JC>caQCLaQeZ(
LPN2Z#UUGR?[g.AETb=BE;<d,\ZRF_(D#.5T3&H+6&I8X&UJP[<;Z-O&UI?a/S-H
9<^&YN^CYeECS/@g/d7QPQJN0g7TbNK/JM2NSXaSGT93&5H.eIFRB16+Y(K2^6^E
82V=K\NZCCRGeP=B=Z11;+bH,=0YGI[N[M>_Z5GMeC;E#R@b]ZP(2],<TV6-/G1I
0aIZ[KT=NGZ8aZIWZ[]+:4D5+3&FE<3=+&WVTH3W#ID<cDd=.+3C9HPFL[CcbXaB
a@dEG6AI65KgO<2#[.7S7^F-SMCBd&cf9@W,4Y)=b2dFDe2?/gJ:IY_7/9E?3e]E
L7;cWXY.@;_>KZ)2bF@#3U5[]^N0\-^#ZT8TF?g7D8SMcc;;=[b=&Ee@O]Q/cYf/
(a]4[345AXWMS^ZU_U68#e6g2WY)<SFY45F2GV]6YQM39L->fEB?&gUXW]#2RV]+
M1cL(Z]@[ON[SAJYF+E&5L:GBCTVG()&)0@?M_N,1Lc2Pg[0SMW?E>9MI3<6GSNc
.f^]UL=I1C057FTH(VHT=.,T./3:LMZM?@J3@[Q^2)Ud5@9+<QP^<+e=E;PF07RG
7X\g5O[dK^NfK3aJHU+PfGbJ3>ASX:MaPNY.Q>;V_Z+_C]99)e4Hae2@RM6_bNI4
Z&_X-5A2a^PYYf[U(/<=83.aSU)(\Re2-=^&;UJe\FZg,ZKP>>Da]@f;P\Qc((f#
?P-UCV_?;)(R/Q.;EBZBP8#b?4+RZCOE)4VfKV;D<+DXS6XY,<;d1FICYIEG>UAc
<;1#LJc[AV3OQ<:SLB=\OA49a41XScd&Z[#,4)[g@>XKNLa3J4aX2X97VAR/T(U+
H\39Ma5AAf15DYW;<=f>=b6_J;D;.^NTQF>fUFJQBf#ceS#->1<3)]_1FL=)L5N5
?Z1Z@1TT[Z7OZ?CD?dYN^_^L+d_YcIPRQF;E69X0L4M8RZDKB;N-KXgEdU&9T:KA
SK0C@=U&P0N9<F;2QP&4<Xf,&&dJYJ,S8TEW9:;=<\VEZ^<1g,V73e#LLKW/T37Z
BaXFG-G</gc@+9\bO&FXDDHONB<>_aCc7a6BeEC0]OF8(YOa6<A4eK68HF+OdG)U
72Cg)KGK]@eI\>?=4+6.>\Yc][DP9fV=^KX=CCgO9.EHP3Y];(4gKH:c0&S-)/U)
?Q]:#WT8KGYQ,:RC=d>R/9/\0&MA\GHG=Jf8#]]]aE?dbA^JX42A_L:MP0dF+0Z7
#P-&1A1=U&2,UX\<E7LD]]DMG829.3)eIA>-/X5UFXH0<B(RX99M(N6TUMJHF9UT
7ECD?.59bHW#C\?OQI\(C46HMO3,>2MS)(E9F_K?,>N#;1Fg-UC.(@3Vd&-YWfb;
.)J>HcL+7&4BN\K.G@UHc54\bRaF\/X?=8H4S02(EXTA(/WCH8:g8Bf;C->QMTAO
E.H;X-W;^5&f@/T-@K7[-OPDAV_C0aK>\G8Egf1YgH56>SA+N3QS&R.UERB[2EX4
PaP316[3-E-/_M^gJ8,)9d;0N.-B?gL@8=@@\TP._XA=CD)M?6/#^1UD<G[9/?A>
.-6)Gc8f>AK(3OM9D4e;+B16<:0(KZ-QK2d&G1E+QRT&K6&F5GFafOSR1eCJLW)d
I4=a^61;/VI11,P.T[TG7TLJG9RHM^8#6Laba>0Y0?O6HFY@T<UN-4FEK;;f12AX
U)D[[R:Z&;R,7<:Q2THAg.RK\[ZdFB&@3G.,GC=?N#78[)E_N)UfUB]g[fB>;]:X
R2^M@<=a0T=dDa),d_dQ92W=[S?J[eeZ)W-+#BdG^[O_XdIB&4S2[L;FFU(=)]_+
>WU,Z\ZK.=FVLF_XS=GaW,YS/#SW=IECE,#RAb.+X=4,Ac,=B]?[3S)df9<(^O[8
-b?E;Fa9b>E//-O7^5+8:G..bcR<JI)OPQ=+(eE34Y9A]2<0(;_YgefVbbbP9Q\6
PeNa@B@,Ne)_^OHB-T^fTG+B@bHEU>EKX/B-,BIBB5gKe.9U/I:AR?X521.E144+
D4&d=B7-c)GcA&J::8DTT.WZIR0a<2K4e8GgHGBR)(3FdbT[7c3:W(YfR:940(F/
fUNdU;V+40LHeE?Y_.5+5JcBBGOK)21A0(0K)e4(cRcPVO:]/<JSWDRNcDVUZS_Y
9+NNMZG>JN8e[G-TU?56MPa.eC.L.CV?c=:))7bYX1@P.-\>FF4C^Qe8f?,,LR)_
/,_FJPAU)g>d6T1,PFO[,ORUCE0=@e;LM24]#EJR:NGV@PQd3E-YUQF+>GG7<\&(
DfX>45g^A397UFY5Rf/3Z409C;aB?8V:DC1EA8=>V)YJRJJR+:Nd48HQ/=L6AYU#
?,UX+A;f9M:UQSFZ,ebU709Z\9Z?+L]ZDZcP,bM(76JV\H^_dI3)[0=L67NaIFf_
YR.@>^?]<5PAEV)d7:c(<])7S.H<-WX^dVa?+3QZcbbT49KfH/@JdUHQ553E5Rd@
YKR3YX_bd4fCD6->0^9:K#@]_&6FPQDQZ>]YVMHI;N3X]NVJ=+6FfQ\0Uea8LA&]
J7dB:I351[SJa#W_U(,_c#M3>DFb2.+/6C[_O:+NWYab3]<5J,X)eR_C.+A689#8
ce^4FPV(F2d.#66VR@\0I_09Q8-?GG59aF5(45X-A,[RF75c(F/ZD^OLa+;EFVX-
>.N:^=HF((VV(EA\5M.0FQ3@+AZS<f+DE.O0^AH=Mb3>Qc^DC67.JeVQQbgZ:A1L
Qd:bXH2BfdG>ab_;S/2J\eRTETYU.A8PAW]B04^V?7O2B/CJb\Y(:G<Gg)H0cG99
N.G/RO&@QRQ/gL@8Wg9?7GR94BX[=Z;^Ze4?>V9)@gG]5KWKM+Z<KP,[\ATfT#7d
8+f1:T0fbO]PY=,SUOH+N:(<O\>-MSYNL=e&N37P-[;ZT22XRH)C+[9dg[c^1UV#
W.X\D/WcG^?M[\4W.JJTM6^d+DDO]2ZWOQD(^CH_O[RC#;Y0_)CR>OR3@g1Kf1R&
_4[QO.ID1>;4:a2\SQ_KI/LT?C7e7F7KRHHW&WRG:gXO4aVQ91E4;7\+?:G/fbXb
YW008]bALQRG2f;E5ISAR138&6^@8E]JDg+)S^QOYSaCP33eXZMVd3fEdDVXb=6[
\Og3]acJY?&KQ6N6(GIeJ0:M=QXJ[?JQ]gRCBUZ9T@E#7<\2=X]_I)/=731+gT&c
S9gH2(+;9:J.O&K0.[c@DG]45^+)B=,V&[<dYL(V.B5gOfRA;A3gX=e68I>-],:K
AY3W-C0Vc&QcA>:EQ,4)G;B[>=5?&^#Q8=K?-^W9SafM1b6dQG7b6YZQ98>\,&a+
0?5f8]BMG8Z_Sf]b[N1&+)NIM>A5/eV^fKD0>aQ?eCF^M&-Ga)-Q&=-KdNf:#8Y7
:HBLSR=P8>I_IQ->21PdD)N47.1fe@[N(bO&]gFOZ^Rb-XA&>G+LX0a^R4S6LLe6
+\+UWTL_?H6)[a&b=dDKU]HGRg0<^PRNbTSP5F40bA=C^/,5T4^.Tg14Na^Q4,[.
e2bBc=31_H5b^TTMWFQHYR-T2-EHgQG/,_J<10WE(c@@HMXDKE.IH>)bHDQRRU:)
&WGdV=<)OZe6Ke8J[O@J8.H+EcTd]H<>SKag\FgOK1T-BBPcGWLNce9RbFH[<W-T
Wf.;\fd=M0)^WN]V&JA#N3B1XY8Wa:<NIZJ<8TebN(OJd;(ITABK)ffT#DE,gNf#
H@aGDER^bJ2:^8BbHgc&YQcNU97\?WML?-XS?B/5SY:W-;RV.Q[&XgRb<b+:>PT8
7I81Ab=CG3Uf##]VGddP?D?&&YgN5Bg)JGWWb9#?cM0U/B.[&8Y[DV+ZOb@cK0J,
bC]TBd-NTESD(HM8SJfg5#^B9Fc2d/gQcS,&G8\.)8-HY]Q][,IU;I-R2IbO?Tde
.TMf_P]M&XU=F9>GaGU)IUMP/G3?5AgH?W;QF#5/SYHO#ZO(V.NX7MEgFUDT?B^=
VT:@F))8B#@@Y=f(ZH9+)0&<V,7B1B6_+K>d\<U797PNU^7a=S>_T=gS2R@1@B(C
\QT>22+(J5/-N,,[IZ:VO_4?7gI>W-N<MdT7SI:.#P-\JP9&)#1RTgNcFQZ]Yc+9
?aY(eD=11)GZ6?P\@WP?.KOA71b_]Z.<(5Zg&+B4KKeM:\E\[:)=Y@J;@ET?Cg#]
KK4+MJE_FcPSe\:S5@c1@eFeLK;PJ[QN>c,NPf@2A<8Gd:C?)4+>KAPKgKcCXbcS
b.Q@1,M9]VRA-:P)TO<b;VRDU<)JL\bfUR^(6B][M\.WU1_S(d<8FEC>;KWYD&YN
V@H,0aX)NCHPT2D=DYL^7a?,#.)g)UXb1O3\]O7>]#8eT7^K&.g3V8_?IK\#=O(M
gQ#B_JeI=KG)S(P_65dF+XBO[5T;P:-aN7TTeB<EbDU/,d7CWf^&3@6fNfNM(<?b
>&?fW#T5(I/JMcOc3X\CP:F^gRW5/2-F9ERd]R.K9/8H[U.eOc+BEG?[MD0@[XQ^
IOVWG^bSU-FY[)a(J;</X@U0cP+dbOAdKYZV=VV+4>UNB0AbO)7GCBQ=^^^FX=>N
1fc8UY<.+(DccG\#BN_Xd>>9_-3<7LYP4:5#UAF?Q[;8Y1;-K/CV&f]_OLbebCMZ
e/T/FU6MKT3H)>#1LH>>,W6#=(Z\^?P/#^J(B6f30&6BQF<-bc/RRE>W>L.dJIRQ
8+R.K(@f9\(J2N\Z1LLT^PH;7K/BgYS9]Y@I^5X:?_C;Q&7G?Q2IO(W-bC>I;CJ3
=_&8MHY];M\F,0SI2cF<MHa4RLBL5;c,#]+6/_>\WX6;.^e)7IfRb&ZF]E3<;,6W
CA;N>;B#=R9>S0a#KAR7gBH^9D&7_&4;\A7C[@fH6<_@YcZ_e_W2^UadcA+Ve;TD
9JL(V&PJ>,.4-TNdbJQ24EcVY:MAM[B=ZZ;XIcg_P]R2SU@9YP&Y:TEdVL,<@[TT
DLVPT5T\@Z9+c>egOUcG<##cHdbS0EUcHF\f:F50_>3P=:0\^/QXMPX()LbA1,+@
fZMTY.1K_P^=6S,4d4I:D,Z,-:1b(IKTG0=N9F\0@=L,+CYYHcL8V,RH\(@g:[8b
=#IY(85_NN8;=^I>GV#Pe-WVBWW-Y@DF#&W]D#f)5:g1[DMKdI6_X)V+NB4Eb\#N
40OAR98-7&5]C/B29C]U^Y2?:>E)dM:c8\@.;-c-=W(/Z?6R(5[_YcZX_1S)?]8>
d,HD?c087K/VVbZ&DU5e[W+,ZSLB[8CGKCZ,H^X?R4,=<?6^5c.\#8?H:We]#S[^
;Yd;FeC@Ke,E<>.<S](HbP3QA8>;VF=2(CLX8#8OL-,\<4<:MB7H>UD<bdJWYT=I
8=BX8+E+,d=B=/<S+CRW+&IY,&@[GIGb=@dF0(S&C)),d+S.?0?KH:DR.BHcWeeK
D/8T@F[ZM[MAA5f3)H;.\C7V<\:^.:)0G4DP<ODA-\<[BC[&+EE_#TN-JJ3(R44?
.A0+4H=d\4S@.]64eI:12JQY=\AS2RPFTO,0OY0^4bE(MSCUa(>&^Q:0S5QaT.S#
31RX4H3/c874R&]2O&G38XX>KLYLT\,RKI.HfRF+TeJ2,[)?=^L-aG2+a&>&3a?4
g_-4W>HT:gP(+@B03E6AX612<Kb_Z?2&5c^a;Z60f_J3/DVPK(a8Jf\L8:<3V]bY
#.1MVL1bT?QF\gP^^[0CIV_@0CeCU.LJ;L#FK2R-?+>-^(4(_9=&EgRVV_/YM,7&
@DK-6[YX8T,:?,CSZeU[@>D->/@@A.&d<_7OOb(fCS&A=)J<GG#UHa6E=ERa>9F+
Y,/f8[K/4-TgD^3a6E1#WG_0JXF:_R.HAJZW,3_JS2QJ,]bXF4(Q<+DSc8e(-\]7
OP#^U+=6c)-fZa)OYIY&LbBJ3aBX7O+4M^&UCe(/b;3UbK?1M-T(+LOdFee1E=;)
JF)_[)L+^:P@E9]6+<g6VCFbPdY?L;Q\eHX-]Y+NLE26C_IcWVNeecZWZK?5P&Sb
Y?:1Mg&&I2N;=E;K]/-M[?M=R)?gG:4CeU0.7.^?:<X+S4W]QK..CSfGaK=fDDRR
_0U@B1@d90dbX-BP;)Z0(7<M@3Z,[TaBIc^\\@+?X<P:?X#5?W()K<[9ef_A)W-?
gX.#?K_a908=45LECfJ^]#=,7S_D1W:EYI;UZ-S9VNE\ZC9_#)IP_S)1e<WW^,9P
Q4OF#8a<=BWFUBE[\>J#4ScUE\4J87\&N^YfZ/aRcR8[U_^DKY;]YV907&NR[I(Y
.07(FDCRU0V5a;[>CR]U;C&W]/]:&&.JEL;]/\3,19<c0@IUa<aOM\_?GK9?9(?Y
I;55RIL48cQVHUZOH88;W]5GSOY:[,08-M+;NOGAF2J9A>)Ec1/T3#]A6Z3;4UI/
98U(Y6C6O\cPLGZ.\?=O9#VgMG^Sa0ALYV]_#Ug/Q>Z/GK7Q+7X3a5g8\D1cfYIV
8K;J>C^P;D)JK-A]HH>[XN692Y+dI]O;02DR0fO0;5&.R/gDXT/LO[_-1e(>OMS3
eYC;See]/Q1>1NWK+_RA&T(H8AdH:=C_7U64DWZga,ba5KIS5FCZ37HS+^\N5H7C
\TBMDQ[Q@>Yc_:+6bXc^RU\B?9W1;L:H=\_FNHf9?M;b;7TH0M?F2VZe.RVIYS@Y
N=gZg6?a1;9UPYIAH<0Sc;W,,Sd]AK9^dN0UFT6A^S)-3<;-)N_DD4B4Oe4QH//Z
^#1BcN?7;MX(YOd(2.3-SAJe.6/IEG4OR;,&KK^0SZO.\KKAL1DX[[F>L,Y<RgGV
2RWMe@LgFg^#.ADXVcTES6QQTJ-#d;b6YG7EEXG:3P#GfA&XbAcOZT<5LSaF<0:>
93D1bL(]RR>QC68NA))HYLYENDR(c4a(XEWY0;H?HE936EUFd<&X;7DO8KE=N:>0
.D=98#/H7GDe5JR&\_>J;7VP+_DFQ?6DJ9dJ;NS0:&F.c2</YLH2H;#PEb@HeE6S
c.AXI=SQ[c\Z<\V@RKg6N@GBf;H92(ZPd0->8>YgQL(#8.6Y=;<RD>e57R309X&6
ZUNFe-2#;V1XQIUCBDEWHK+H]JS.,5.(Q1?.@<d)6(ENMC:2G^c)MVW0BI<<NW9-
)^VLWXWQ8IJ\81)VM0M@,;5=]_Q,f[FSW8d0a?_Cc6\79e+55URFY:P9BGEJI+LJ
QDEgUUI3778c\.4KPD&_\MLH/gMIJS1G_cK0>eaJ^L@H;/>C)?X2&XUNW4V0B]@I
U[RFcZ?40a-8^5?^@?FK?WR<2P>2)X90)-&0=ZH3YCDN#YME/_0J-X89DL;IJLQ,
A&V+5T5;?d-R30]??N(gCg,0+f+c6B0,0.T(Q&-0aVVR_(>53?09P>>bQ\F:a6)N
g9-I&b,HAC&YD@VSJNbQ]<f8(-8DXd3RA=C&=OUHc0+/2c=E2696Q]BUTRK):C/#
O^742]fDC_.g/>^f^].P,<J+K\@<e-X24QP9@cDCaP>^5&QCILaLS,4_FQQNEfbe
/_D[<bEVb:EW1&3#>bR#7Fa,Z81U(^GWJ>@-H]_\\B.GV/JWg3I<XV8N9/>Y;=g@
6:YAZg>^0T(Y#\H3dSE&Oa2+/=#/,O(E=0VHT=W26>W,N>)3]#7d9LXdH>0><SZ/
\a]bD7UWe4J#\P@1d7J9J2VN1V6YZI_aA0KS6T_#+G4,b45N#S;DB(:C/[1U340E
6eAC4>bf41V^5<]+TX,W7#ON6AS7dg3SMN)V7ANW4g/4ecbWf>Y)N25_N0^Q.ND\
-fc/ad+e9eV\cE+2C:26cB@L&LQ3LFLP:D/SdIa\ED-N5_.S.7NGBX[]6VHM6EJ0
4IVe(e)?,g&#U/R^SWVD)]U\<@LTJ-OT5/.D&Jg^;]SR?\[dg6Y.7dg7#?,>MAT6
8_._-fZ._EQ_9TZMF6f)=C^XQ7O2Q/XMX9#Kc9+R9<H.N(M7A(8M&+1[c4;:1]&7
Zf1gGI67,\^L\7<03E.RI5UC5LZ9&AT-F-6<ZI2B1<^TRI>QJgB-4>\48GUbFGdN
?^X.93bC^>/VER?J^:)3)94,/:WNH+E7BJ[.&XBX)<^^#F;EVLU<b3;(@DG#1N<S
Z67EVI8:7WN8dY?H^]:S#+^7+;PE&I45JZR,FATODbM+B^J+<0^f)@CYE?1ceF@#
=bgQ(ATGXRQSY1b.F7GIBbVGHd?.4G.\2g;YNW4)C3W@)^KV7^Y?fW,_e/.AOI1d
3=S8HMA<[6E/Kb)T\7&f<92RD<b?c^]2[,Nc?I(HIT]f\1RBa/4BFI-eK0..8H_O
fOgE5BN#].Y0,U,Z9>aX,#L>-^N/7H1c>;Z)c[<_>1LUQL5(P6G;7>/9JePC)MH4
,9M]L<=\.VI?Ib4[:0VXT.B?KIML63<RL\U+\g0A.XWJf(?\]_(_ZJF;U:CU3.2\
H.RIN.LRNI+9+a+NE@0.UD@5U^7V1D#b7T0,VQ__+d#9<J/fDCA2.3Fg2_UB+8+F
=V1,UWE,DP>KKD-7-ScI0I9\H)U/Cg[_S?:f#B0&<K^1/Rg\Y#c(^Ud47G/eXcbU
]8.c5?=0PL,7BP=P2W#cb9:T+1)],AVT?CZ6Q=2(6gL;@&YP56T;5(H>L4<V&7B^
)Y^O4#5ZB5N19?)L-M6HfDU6<ce9U29B;5Z(Pe]I]OZ1(RdE:He@])OM_B:=C_.0
c62N=W=52W>AHLV.XefS_NZZF=Cf,5U-EE]a\-?U^;L?J)_J#R5\G\(O@7-MFOA&
8]K:/7a?A;CR)-M8MDYba)7WFYJ>,5?-3PefN,D\beG6@C/0YX\\HUgD1I3=g(;7
B?VaR=BCVfP+A>HREPEH\e8H\NV=^]K8(\@AN-eOf,K@2e,I&A33.--FdVEHA6\4
H@c:KTLV6C80EX&G,2:WJVd.ZBV.KVB@Ad1Z&]\(AIJOS1eYVR4>F>WJ8<S?fP25
gUTL/X@EQIOR/<Jg5Tg-86TTP7PA^<>=CJAU?Yac4F;(;Jd/M]dZU;PgX,]+00RO
Y]C?+,,4b^gX5=BI.\3^f>Hg.:Z5CC^L^[ce3>DV_D4V9_D^MG]WWC.dF[&I)gLO
WNB7G^<Fc&_+EEe1JdN&93,1GMM7(3gf@T)IHOLVC/#/0<,TOWB@H53Q_^5;gGgf
H-]BfCK=HBUG59DPI85Z([+6AaOR5-7H6?IC:=(L\3W5GR;.E)N?70C&dH>,S:H<
/=R8UXJ0&9=F#D6V&=YD#KHAMPX&#NgSB\Y2NC>?4KB]^Z+NN8TAELY2K,g4.:M[
CIYScJX\Vf=Pg+bA:)Mc.^UW&=_26/CR//-FK1LeLV/QWd1&^]AgY]g7R3JH7W1.
G(4a,C>1TYdHA6D2N>PXV+W<X=A.JPC?AU23aJAc#Y0I90-9c55\a_R#29.7Y.>4
Ka0b\=62MQM,\SD-YEV#f@,F09;5Wb6,JeYYETc?Z2A6I7#TXWIFA<]JNES)95;2
5M4_/__9E+)fRC?RK14Tf4aBG>6JQOD=PLD+OdMV(_-O=VCB83eEK[7YF7cC)@6H
+:WCBTO13ZZ46A;.Q7MYB9:1L]?DRa1,NQAR6B85c-X,RVOgS)-f(]ggHJK#^J65
E1gB<GTA.Wg]P^gKFD4MUPTV87&TRDI0f#;_gGJ5P9e4;=PC3S_//J4:[5g<]TIb
GT8Z2LdIR:,6P>7^=<eI&6@_KB4?&Q7RO]EAd]eE,cF)69W(b=BXBg-fB17MU=4V
]cO)b3>M+-WUE;ddD[;;G3b,g9MOW2<2>9\?ZR;Y/;RH2TI\V1Z]W\,bR3bL3d(R
M0/VDU2D6>\;G^2E;^?C;C(ee,OQf0:7JF)TV(fB[>a8O1Uc72=ORVMYOYV\e(ZQ
3e:H.6V0c>Kd9L<10c3MA5I?#=]^UH=F,);N1]d_NJaND:;XB8E(W>(_VQU7@-#K
HP([I00Ed)Mf9^cQe<X,RA?MP=/)E7H#VU)Z4TL@D,(TX>2g&2NL6=T[V1GF\g#a
Y2T-87;8:[a4@]N,J\\/Ha68]GD/F85]FG9\&]Ce0bGP:0cF_dU;V]Z:0@/548VR
8C6)^\&10J9L?_?QENOL==:8@J:-L?8dS_<+H=K(cC4NA4/JG<G^DC,:KJSD^-2D
f.HDfdXZcKPf]_5<X2<@VXOe>-,J>Hb1S(3WgK0FXU2H9):P6WQ01^5HNQG4S5TU
V^AQg.e^Ccb;PFOfEL-R[^#K>Z;N]CY,.13E7XGS/7X6f;FH<H>>LdI2E@5G8SA@
9AZ/Y[\e1J?=2]V<75=:WIMD-c++D\EMKDAH.EAZ_C+J5LL,TbS59=8,b2M<M2L8
)THfY.?;BTb\I7PYf#(>V]4RP+P.4JB6##)=cdB5[H@W>[;H=M(P2\K/\7P>Z,0O
OTCL)<JE[N)IPI:LDQ)P;7O:UXA7M8BXVO[B7Jf7/#7^a]QF<)2Z@N8=cHDKZ#]d
\aG)Z0:XaQ.df#=[\Ld<Q@K:CJM\.Z9?O9SUVc0A<H]1,fN,@8D34PT5V6G_>ENY
>XV:3BD.;3X<aSFK7U;+&8dRUC^,D8V]<g11E[b>G@=#+_dQa(M2-eSDR5Ae#KJ+
eKgH@;cbbSJ[3[_=>HXIF.+8FbPD<9;X4,M^:GN3]d.XZ^d54OC]#:X_5B0Y=0T)
fS4\5gFCHNE+^(=O+J+O/P:?(2D6TCN,I=E8dWJW[SKZ;Dfb@NGGOaCMbLSbAF1/
WIZ;&d:CSe3J&894LfLbK&,NTU\KdH\;V-Cg?(3+)dRc\81R/<TGD_A.]^+K5=+G
g,9/0G((4X^b(U_1A@.#<eIOUA:>#g/a1:][UAK];1+^F=23.I0CSR>97>A-^L>&
g74DHO,N<8ZfeY?4a+&&V=M<UU7)X1?(SY6??MO9Q=cf1X@^UL4X5dbVXf\C<=]G
C_#3P]P/9J-FT+<065B:5^L&A0R=V&J90@6f\Q6MEZOA@([3N/4??4dO+#RM[(?&
b,4O/JIPL##U;^@BGf:H>eV74>@IR2,ST2+2e<680[2[.dY:^V@);]AIc(DJceQ_
_X9&KgBf,L&]HU?<WQP[:PGE7EHc>;A7f8[1cU:fQ6N)57)U&#W.4&9fHF?GUG85
;0_G:CV>>#I@P/,b_,P.F5-;ZfJ#a-8Q0Q(a;9fK?_:09;.N8</Y:0e+?;P-<>TR
)PXI2=U(EQ<X:HgA?//.;I8K27C;QAD:WgZVMFbJ9+c,<5W=)VeUGT(1F+^JRO7:
E<>S2F<_3IJWL:]#<>68PT8Q<Q>09SV1TQQ8bMW2+:e]3QY\K3UWT#N&3D@aYU__
:+P89[9RWdPe@0>9,LQ3DD:B>?g^aLfaB5WW;-&BXHR5cdHS+^2P49(P)]95Q(B;
T>.)G(XKFG[g4eG^EQKF5H;(0D@8V#9a=;JT]E1PS#DYW32FeaDQ5KW;T;(,J3#W
>2JK\2c?eSX+:PgX/GH_G^:=JS@.VO19EF=3R96H<.-J+Yd)&#cB4WUB8)+d#ZF6
#:[8B,F/(R&3QTC((-;SPg_T_cEQ0?-8<6K)UQC>LT]V3X;8g4H#WO\?g^bHJR&E
6EZOQ>.CeDC\ae@dQEI=J^fMQI,TYd1QbAC6W7L^bYVgJ[e5>^7BJc)X2cX-F7g1
QE3TJT_:N2BAE/g_/bN?cJ>4Y69#^X@(Q8gYLI+a6GME^5;GG,9LS>d[@O(607Kb
:RT1O;<[-[6^Y2eLV.?5^PH,1G>L8V]fb>B#;UEgK--Bc[@1CY9C&>-YOAH6Y6O:
dMB6YFQ\A7JHFO6gW(@UCRYO0V<\E05FB03J].I(.I6L\#Y:[BfPE[MPa;,,+8]G
PW/>W8D.3)A<V<d7dfV>=@XRH&NL(;WM<MF,+gD@VN?#:9?d(F](Pg+JW,/Y7gD-
7\\f4C5O^Q?H#;W=(AfPQLU>?M?K<.#-9:,.cC??SN#GHdY<D/A>)?;\&T;5K-<)
f>eX[M:ERY12L(,]ZE5S[3_6-c/QXHSJ#N0P1b&<9([b#_]V8f(,<MCgJHgF8#PV
J1-XGfVM\D)[C@SW;<(Se]T+\L)32U>?YE>KI?SCdMIG,0:&(>0REgX_QE]<#e83
A;Eg9[be53+N&0Z(@POC,J\ZS,D.<+CA;f-KC9Y&;L&G[C2]fJXQNA&X5e^G>>Oc
F8VV0@0^4Q@>13]T1L@G]aYXAM.f/ROHd<<5NIZMS]c&<:I/ePD>#fW8S#).=:+S
J<93>\d<3fWZ#<6A(,Of\O.Ofb+]e-dVE5W8/8RK&Z;V?PB._MW(>_eD1[V^E/_W
K_NHg<WD6.,7f,K+S4PG(R>4DLcY=#FOVF4U&f:;TVQ04[d4L8A>bDEbF4Q7E;?7
Pc?=_?M[-8>@J)QJ-9N9]EXY7ZI=8HV<YMO7RG7-@TabZ,7e_D(Q?C4WHQ@B>Ya+
WWW(;+0V8P0:dPTDQI?[87cKPW8&7Z2&6LBYEfQ&YDMVcF3U>;2Q:AP+PKXQ\O<U
D,8M7[K@<aY>VP+<GFCagbeB-((TI3Cc^I7,37\3[KaA\FIH,(S0-0-TBX2LWZ\K
CNIdG;UO_f(X[9bFPLM09I^N?=@g0KPe=MD=#I]-[ENQXbYEE/&G/g7)XNR(/ag0
U(]1g,cS+eQQ_1\G7<;bBM95Z_,)N(U.09,bG=&);LJ,A(/2)FV;-V3eLNT=8^CA
8ES.3>#<gU#ST?ff0LSQRDU?594^5a8E=BG)b?KI\KBS-VR<Z)7OXVG3]-a5ASE.
=S<@;L)-PdWQ3[Lb1NK^a>.]B=Z/Wg(V?81I&.,.f1F@.@CO_Ka=8,K]YOc>4M@U
Rd&f9HQ/87;^S:[6)ZB28_-Q+2Q@\DNLEg(@.7GYH]9W:OA8;Z1?bX9JOW=OV9=V
<+1,_.,;2S.FV8M1,6HZI0M?\Na<P@b4M3V:_cYg7+gO3?E6Q,Cf>4Y;LLJXWKVS
L8G^MS]BP,^.-3b)\)0C&LTKA5(/<D+R0fW78Ad[dGHKZ[cGD9dF&YgAVNG,O56,
<T,a\^AO>dUIDa7/b4,GXeM+&:KC7)Z__J;H_b\Z>e4-#_H5CG8\6b@HB^B]4SA+
>8Ne/5aM)3dNH\Md@G7(&9S&-UaECM)7d37^>+389XXGD8UV03b.ME^TU_#KAbOH
:.1HXLAMX_+_(M)P/4I_SUE;a>R9OG.fF]OEC.Q&91g.FA(MIJ25/N0DH>#9L<,I
SKc[2U\#NgYe.W2R9C5;J-f:V+H)TdEIGZN@]?1)H6W^6Ja#[916S##0C8#X3)Q3
6A([4&D9,F:XP.?KF=N-93QI/U18CFI4AIB7#b5(F-@ZDH_HBTebYP2_4:7,]R4C
WXK-=gQ5==WM)aS^:)&\<b3<CA_E]Z^NX[_-L^ceS+[NRVbL:<S[eRWY,[&]6a:[
4f87DYMgHP.1\5M,00G1D;9.LaH\K&f@^5,2]+.#]2Y<N4.YC^6UQ3L]9HES_F=.
H:CS7EBA,f#baV;M72O1N.@<(Tc.K408>B<J<>fP_<C1+#9OFQG\K6ASBG11A[Xf
V^g#@7,6A/a=3Qe.5#O<:?X94Da(YRQUf8+G^NY5J)F48@.IJF\>QQ(M8.5-13]G
M/A?G(L8HH624VMZc<@Q.540E[GT/#).(B4B,]UIDELdf;A_XM@R:@,=ATB&dE=N
SH[II-cRU77cVJ?,[-TDFQ@8U@T0L?8c[J=3M4-X&48Q:F(5TdIS\P,NI2);RMOe
+3+GKEV+N3c?/4V&[#Ed)bG7)@KY8:Q+3/#FEG#U70^HL09F+48M47)3cX3(Z[Q[
f4eWBg[,2008(0R@B/_/B45J]\aKZ4]:>8;S9&O_LWd^37#X1J-IM6/=F+9RVZ&@
NV[(21/ZG<FafKMRWN\UX81d]I.]CI.0T?b]&,-H_6L&2#g:ag8#^PVVcg1eQ[b_
4\B5EHBUI#@ZVV8V#M:VQ,Ic(K4<4YA2E?V6=7c[F#M)D?A^6.3+?W/[ED5CYe]]
2e#c87(e<U<eGcYf8:RcC\ICe.-a5F5-Q6R=Y/YL1)P^^G4?fcPeG+Fa_/-PYU1P
4Hb-gLb,6&:DS9?UBH55/7IR[S/0CJ3\d<O_U1<_-JN#0a>8+&3&5ca?cT?BaU.B
dW,U?PR#)>d)VP_f)>/]Ea)ME+9:3Z^b]QfGP),U24VZWZ6E?]=+/;F9D4?Y4eM<
JPB?A9#b?\<NbUcC(Ag.#92PK[W<TUg8D<)]4H#>39&D&?c7a3;g=fKF4E)OTG^?
6QM307M&&aMFV1=6V\c3]ENE4Q9Ge-<-fA)DdDSJYO;]5;0_P6S-<AORgc/I/4#?
169LaNdG+HN;7N36]5gJ#:Xa\HDe.TOP6eQR?GSI]^?LfOg\<;+9<e>^3bZ259M0
^B:bN@(S_<@;/$
`endprotected
