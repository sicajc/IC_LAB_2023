//############################################################################
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//   (C) Copyright Laboratory System Integration and Silicon Implementation
//   All Right Reserved
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   2023 ICLAB Fall Course
//   Lab03      : BRIDGE
//   Author     : Ting-Yu Chang
//                
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   File Name   : pseudo_SD.v
//   Module Name : pseudo_SD
//   Release version : v1.0 (Release Date: Sep-2023)
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//############################################################################

module pseudo_SD (
    clk,
    MOSI,
    MISO
);

input clk;
input MOSI;
output reg MISO;

`protected
H2cP&AcXK>[>G5GV=L#R?UY(;(24Qc@(dQMeVT?^_YR?7V(&R23:))EV52gME\T>
YAMYJCe#YU/72:RE0)f(CVV2DP[I\GYQ(dIgE)?1G1V.5\&gdI9W<9<R2fFEH#S,
B?/I#dEY)1)?:<MCbYY.Jd:D,e7GfM-<[<2b(.1?&?cHc4K3fB=Z5+Id,T6cf>g>
\L;<XN@^c=FG\a(8HF\OV)<D4JZ#=3bU:HU_f>F6=d<FE-^f_UWG@AW]C]H0[:fE
;3,5(1#_e7ec18V]^cW43?/HW9TCXVMKLQ:PUbH2/9[ST.ET/.TR/.c:P#7]dDZ9
[@B-U2OF)8WUdA&/a#Q6]_KP?44d&79JATON6D85=+)CDHV/IRc@+27HLF/Y>Le@
?=M<1SYS>K/@[5]WX1K?QMYZA2FX@]LGROJJB<Y(25?ePA/gC+6]?H4DC<2f3?S:
cFb;E\G#FR+6[51O_Q?;\cKQ>3ZXR?RPKL<.dW;<VB-AIE3]EH=H/M^UNQ>bO#Ub
Q_LeAb>S7U1MPQUPG6W=L[4Z:UbADV,FES^\>9EbRUgJ2U]cABR(;=Ye8-6gc1=c
)aVU+#@[?.+_AX8a0TD?<\W?gZ3?NX_>.JN[?N]XSff]GRK7IEM]DK&7VZ8R1:7b
UYD0f?M/5Q#:aT+VIgDI1CG.[GTRNE#;-e>eUIV0M0715E[I\2?bR,:gc/I<[c];
eM:^>#G0/ccG1QY4MWg&7O>:\#c5DHKM5-_I.V:EH>L7#BT2H)&AJ#LcXUC#Z;27
Y);^#7(#eYK+<0-6;NE]F@1Y2fOA2&&0=>HT[IDZ+dL&9J3+^aS:F\P<:B#>TcLV
0#S,RZag0V>[cPC^)[__QWbJ=aV29X@de4^0<g#HR)F=Bc>+3A;Dd,C[gD13WW[V
>Off3>T(KMNT2X[EGA92]SU2P_23BD2@T(WRKd/P@OdZQ[B(TZRYWYMeX_L(DFUY
b7O6bfTTS6TD^LJU;P5MVg2]Kb0QLg_@X9^HINF89-EMZ@LUUHV7Zda7:eYc@/g2
E]</HB^X&4T&d1/,:;[[.I=ZM#6>>C_6.WF=@fSX>1[I5R\P?-Hf/]W2cH1+R4A5
LCFOZ&Ua]9.XX.@02^:3VC-AfAK7g@UVfSLC69E6@?\d>g\<G9U2A@aS1-N^,&-?
QdFc>Hece2Q8<;9Yg?_N4@c;+#BP\,<a4O2dM0(b-3R@J]D&H:HAHZVQJ+R)71,6
G0]S.O2S<T@I:Lg4J3>X^ca@2=HRg^O^e?9UPAgfDMIC^#QRU7Y7Ca^Q(X/^?M/L
[Gf:XV9(5:F^.c9568TCdFW>8FU_K(HF-8KIe1O_<YKd8C_C-E-?(g.)WLfAJC5a
[Pf0Y2.\8ZCIC8O#dD<X/3UNc\>JD#0GL/M<UN=ZPT-M.[RGY>Xd^I;@?K^eLA?R
X34YZVKPSCX5_OOO=\]Y&1(ScT0,F.fF5b?VH@)?aL#_YW#2);I]X56IK0:WA?W&
@53O)Q.\SbNUF0O9KL5NCLY/:-8==+=e47N_d>>7QfPa:CV\a)DZI+8CV>QY+TVC
Q9CQc;<f;9.;^#?<XBI_FZZI<Z(:@TLb,_QH6K9RaX]CK+)gPXdU4e,U[9=,&@BG
EROQBa(?Se6QEL;8ZP\X+NOK<>W6]X#5W>c,2ST-WP\929MD;Z0-+^MTMA+,^IGf
U,fO./&UFDg1Oc\b(.bDUX;&6Q\S2b;X,77N/d\eQJ>T21[Z6(Hg@K5B<BA7VR##
/EaZS,D^3CfH;4f&&S,34;V><g6/;>TV-1H/>dfY?8QKW^c<;IU_c[_?1];.L?G+
T<JGNFB_T4?PNE=HE=._fe-,0AdJM?OHJZcF)-#]>IZFU1SeRYZ>1I:/&EaeHJ(O
59+52f3eg+@da)fGT<1_2aH/-3+?#;+S)BU?0=(LDC.D&2f4Bf=5M2@&6bN20/-S
)&_D=KM5W&^W]d&Wa1U6)H13TI@LHfEfVZ3c;@_8^+)HYcfS]GM0&>&Z8g4+US+f
RTG#f@&OB8&-H]?R4&^_eOM2UYdH.,^N/;a^[1^XM>fGg7R<Rd(WSaf\Y&=D2/J\
?\_d<eNLL/BRZBY+Q[57)41L32L#+J#_Z-PSPU-B)g)NRc(/O986-Ggg=bST<Td9
T^0)bF).cd?BFXb?+1@_H4>G?,AV51EYT-7[(]aR?[dG@DI8=R]G>YV#,HeWKJV^
PL&Mf;YS=Lf2?14N]+LB&D+D([4PbG:R,16c3^>ST]R)=\E5a7f#?//:QH7.3;Z/
YRRGOMK+_0SaTE;N/?:O6aUc,&WU=?1TNZca&4NN8F51&K^,VPZ[5dLS68+]8\/4
I&bM9JUcP2A)H@<4&>a,G;QRDg+Fe6H[UYJ;K>U\OLCXg@Z=T;TbEAY_L:FZM1S[
3J#Q_b]f-_&2A(cQS^>(_L=WYG_HB()<F)D35N_>5L2GF&-=<ZXNG5e,BPYBAgF;
;aU7<L+[cbH\KPS2fU]eSET[JXL&[R/6PO[a+&EC<Z.8WXD<6HH>cNL&#U_?(ULg
^JZ-[OJR_@06RX]HN7.HM;4..L13g&Z\)F/68W[71?D7OG7C9MYXfJQgeJe3J]T4
\Y5I;M9eTMS?)c[73[HDL52[7-2##1_FN(C0PP31:3T2FCb#GJ4SJ79O\ba&FL78
e4EcE^]CWP\;aM#(Xfb>70e2NPCf/ab]&KJFYd8O/WL&5:1(:RV4Ba\^E>(4WT,C
K42=::-1-DG?JI+97HcU6,a&VL.+L4+X_#Mf6E5fQJ&PO^=/2DPJ->&Z8Q03CNFF
_acJ[9&J(aVQ)L2g]I:JCD:B@8^2AXK-;/G8O)8R7\@A92e>b<K6VP)W61WS@B>+
QQ(W&gSHWRIATSc@Y(L-3eVZg[S0L4,RB]6Wf[;F.<A?4Z9>;C5M[Y7NH)HYP8Z3
=.f:H5gaF/c>H.0_fM2fB<A859W6=XRXaPBP4A1Jg0)faM+FDf5B\8O#6cd)J##)
;D0KNV4CKW-Q7+cJH/P1A4@Oc0:cO&O:I>d<&-(F.\<3A-UA3DAdDb-#TT7/OGBV
1FJM&NXeE5TOa53.^XbZ[7?I@8A7aH4QW&4-g>?/K;>5BO?7&)=HVS(0(I,RX;)?
2LKZa[^I-Y0573PR=K59P\;@=g/=E&JNMaQ?DWb5RM]OVg]?DS1ERK+=8LGOY<;Q
8:\7JTg<<ca2.)5QP656a7NWOgd]R3YX;A-cI>df>d3C1_^SaK72I@Z.G,FI;[]N
H7JcB<fH?LcdZg=40]ISVM>Jd9_+]OE_^DP9&S6a&cg7LcC2??cBF>H_CWTTaVJ]
CaEX3Uf7S6NP\MBg.K,TAYgfdaAEO[.B?;B1.N+9g+0:T:c=S(GEfQ-M^@PC]5bG
Sg5B0/Nb(-6]J85DP]2-TNXK\&d8\XL?T)2?<X-DEK@7Dc(5;WGT6-QAI;>1X:#R
#5=M[1U&aM<.+,YXH>SM1G5cN>W/Rg]dc)U&b_A1MgW@_V(0F((\GVH2@Cg-B>VH
C96aIA0QPUV@(aQ1)2DI,[Z).&dgW_W\R+#M6T8c>LS6<.+ce(@C.P0D[Qa[&3;e
3f0d^aI1eCAgL@<G[c<-R-cD()Kb,AbI4V3D;+IaVGYQdRO<?J@ga:5Cb6&b.9Kf
+I)dS[.g5<5HeAfX;M3F:=.X11J9D\W2./-ES\I@[]]e/EQJ<QF-3L#7(b^][MVa
:/^W;19;WIPET>H[+<THfET9\/ZQ5-&fe(/5D]eEE#dMV.#1E#;H8dF\FL3(Z=00
g[5:eF5;Oadac@+b03Rf_A:N0I0F=#S>Na9(S6TS)e9;]_?@LaEf)/AEITTcXYGX
<.GNG,32DUV?C2CRL1>+bW^\,#VBG5K[]&\(6N5NeQZJQD/]-LF).M5DWE&\2ID&
<aX8GcNW2?F5A9AP#[U-83g)^c2GLM8C?BID<G+gce^d-6Q\#;O3[R=0BAB&1(@=
NZ_#==9OWBF@#B2MZBTBA4Q92,W1J]-RJ:@8c)E(b@L/]CTEHJO5>dW2#F^Z^\TP
#_G30Xe[>/&KN:&6:JE^D,T6V_Q=_:0c7&Wb4)O3dAD;6#BZZeQEFG=OT4KP4>F9
(D:+@NDE-2g>V.?&,W77V<;>B#O80a-c>+3;K:<1:A=PFg\HW^);I4URe6?JVDF<
a@^KD1QQNeE>8+_\BZ[9<Vd>&HQ_);BU)c>UBSBD0(ZgET;;cZ;@Yb/JY?9A&.Q?
(g)6>/[OOI+H_+d]+GbQW7@IOSF64\=#32:eR<9DZ=]JU)<WG:S/\,O=dc[Od096
RFcO5I.+Oc\J<60.CI6_;9\-^DHX\Z#590L3@X26R8fENKNBQEde4RJ0QMHPC.P@
X0/Rc+[]0.<Fb\-]4.^OcP0FG)EdeY/L&,U/=VD9Tfg1C&#bM7@bV4QR[CO],<86
(I=13eWdGdM+AVO.IC5eI/e0PN=UcR>b=&UacP>aT\?L,d,Bd?H]:)e:)SaV>^NN
H</I_6FL@-5f&\e-LBQf^1BSP^+EPVU/CUHT;<F-OL877#6b7I7,0?^S^e:88JN[
@UBeDF+&S[)/24^W;e<S-Q6\CKT<?RWF7=01&0[]M@K[9=5XXZXI/D?Ab)UN:.Ka
c&F@/MJa4\MY+]N(f<06bdcG]3,T&GAQg.[TUY@)Qa,=aGRgV5(I9W<H.+1V;2_+
>S@X5cTWQB;V_11;TC5IM<HLL+WQ6N<Z(A5X=UNO;465O>cGN9UAL-NF57V8FU-F
3AZ<f>6D;e>:4QQd-X:#cE\[aO4.>(3[276&/07Y8^9OH?[I#FZ7IN;F7&JQ:X:W
^bG668AXX5T)DFM)b+fXNG=^XZTYbEE@KCVS+]M.;g=5a62b,)FG_G8I@NL4+K-?
R<cR);a2O-<[PB[\XP/17#<GaD4?@);(=F;[X<[HZ#bV?TCP=d(g8FZWAc+16_RT
SYf0=;(#YQA[<g:FfAQ,P0-g51GC-3IdKD=R+Ee+Gb3S8(MLXbaYc>ec+@B^ZEP2
^[YTLC\aQ_f2+BP4<\?O(_(/80e9g5-OE(B8d00D\>,@^/@[BJJ?[U)<c7_7LS.=
<Z9a)b29S7RU4AcD=FNX&LGG[5#8)_bAaF(<K(U[IQ2LR&.>ADg(Y\I27/JU(&cP
#3>QS)=^D8(B?I4Y9-OfV/91TL&J51J\IWZQ8RP+dYL+</_gZ0fPSJ.UW3PK5PN]
W)N20GL/)U[\#W=D)GPS3(V-b1./BY@F?^.c4)&P;X[5A>FY)\28:K#<&]XfR\de
1&4/]0Cc7>]3ALO,U[H?TWaS/J2DE8]OQS>d2TO.:5Z?(8/^S#QKXXB&J_S7[UKC
CfSTOD#=#\OgS:;WMgV4;d-[[P3fC)--(eg6\.cW;[M]<Q(XJQ3:@Rd35NRLUS@4
:U1:S/8RQ<B\:)K+@U..>14QHYaM6B,c:4Wd?TS):1dOB5G?=X+J<+>D?G]Mf=U]
>7]LZ(5bcNDAIga64?6RHe[\]gJQW1W&]V\E2Z^-ZU=+YV>W2)Z.6425U[d>-B>+
UC=UDU22]g-H>:f#C=LK)WEKDT>_@9Ka9fK#X&RcW,Q=PQJS[_?]Qf\X@GZIMHa_
@MI)]\FgN71:SNXeTKf).(+E94@+U?9K+MB,AbB4FYMP;MI2e@R\]V&++CE-CZ3)
KR]6XVMF_HQ3]\71_CYeXWYD9)dHG(e:+a>3;KH@+N7A6NAEG&cFcBfab3fCF2ZY
dE4UdQY,#Z=VcR6/L]6Z=<-3TUEG3R3KDV\Q_f?.B,]U+SWP^X\GGJ0=0D@gMH=:
3PID+UKM;Bc81D(._NL=a?Hc^5fPH22:_4AIWH^_4bPc8g(c6P82[:H[8;]N1fF?
F:W]0gceW4)/CbdXF21\/(LL?UcTfBYKgaW])6ZOBYOLN]XC/JV:R_)K&J9&W>/W
[3?S),&;SJ0>DFK]=:+&.5bK#/:YXa,+/+KQ^VF-15aP^JLUdXFfW:E;YR/J]G@E
_H.O</2<B+8VT^#,^VS;=,LP&eYL7:9/K]2eeF/EbZgNg4dT0fgA8FDIQ<P2G&>C
a3#G2Bf93c-6SUL<>&JC1_QK6[H9E0O]^9&=^3EX2=+DVX)ID>VBR];a+aR2/E4e
E8PPaA)e[(?&1PeaE(e<@?BHZ,L8?78f^7:A87?]@>G1+D=5\G9(LLA?SdQ32F0/
Q#<2aE0=S:M9E3(#.0)0B/1HXC#/W4=W>@_3:TVQ-Ka>(EO^:\MMAb]QUP?JL@Ee
>T,gZcG70T#[)eG__C#181/<UXb[TX0+0S,SJ#P55F3cF+g\eYNYZ5B)^U.ZaIOa
-,==3ZH-FSgLIQ8C1c\fd1KZb?BZ8dOU6H0^=N\3&:THD<KKQHU4b1]P&TcY8cbI
:QN@.52TS+a8DCNSfG;56:UcC]Udc]?/;?gYS),=Z4Z#ROHPF8NU5J8TcU=RU&@Q
[F+QX#)I).70&QfYe:M]W0fC=1L;-T^J@g88)a_:R-UJC]B&KUC(d_;6\fT@H]Fg
4T8c/+g&6<\OAU?8O2gJJdH6Y2R<N.cdKXX0H^c.P2#dg&\/HbTFeeF.d0gQ1[11
eBQe>:H)9?fcE?4CHDLE,gfZR_OT;QA_UN109N;a3B,65]Y.GeB[34b/8S+cSCWN
91ZQ7O0J7,B]e,68245S.B+TM4cSK>(O+c9<QS[-MI;;/2)U<@QIY]VW/SQc;1:F
MI7Sg6Vfgd+#EVSJJScB^]MO1<3>T3G:_g]HE@ZC))SYF2O<)LV(HJ0VE9-/C4aA
Md=YB^S<URFOJReg=cHVPGB=ID=G&fP+;9[&S=EU&9W1D^;#JOHTW2<0bR(+&^(K
(VbF&?LE]6RWa#&<S7?NR;e8G:c<7E9\ee+c@U6\A9<CTM9a,#Z_YT8e?WRc.TJ-
[a@_Me5EIb[C..+][2:(]Ab_7aH1DV9QTYVC37Rb=VF(DfbL=T1Y;E0^X4#b1Tb1
@1ZU&gPHOMQ50VF-?,]De7S0>[\R0P\K\<e;Q8Y4G0/a6Be:-\Q^&^WdXUI6-KBN
KcN=)YeAE63Xeae69a)J5LfTH_HCQ72NSJgWXgRBHU+/8ND/g6g)@O\2JF;;2#V9
d=,VdM8PB[?0(0(gSI;QRB:<\13[OFT<J>/KZN&NdD,H-75C/PNXHEU&&0U._OT4
7[-:PTcJ4-@bZYP&g4IR_A1:VI&cJHBP56H91B)LUBg_eR>L5&GM=N]gM,]U&.a]
c0U\NE69e0b=1A)1PK0@0=7<<10e0V04D;=81^1FC,OL4MFUK3H/U+f^.VdGF5_K
T;@,TS6(YbMR.g9V^-9Bd>47Ea,fMH,f8[(\(HXZT1_dWPSI8D2S(X1a=&[<1##>
:M3#C1gB\66(Ne/E[])K<5H_2/KAQ0^E5S2:e1EY;AP6;L;I]681HI2OE+HY#QAB
=F-D:?Z._]_E?U\XPS5/?0Z/-\T/W;33JcOBAeQ1NAAZK&N_2FXLZ?\=>.K^f)d#
CL0c@c+#;c)GT6MFg2,Q-)?CZFZ<\<;\McE0:5g\aIQG.:YW3UV,5C6fE/L^ECcE
6F;._gC<dDH]G+0Y\M?D;[T.aHJI;Jc.cB+\\1::@,;\E0EQ#H/dg_dVDP;Wa05f
PIX[?(bTc5^]4((>K842JJ,TXf>BM.IMX?85>GOH2,g9Z^XQ<;2<HRXS@_5_C4Lc
Jc.3SPGgRAc;,g;\Hf<58e&f9&CPJ)fPZO.S,M>E#5M:6-@T_CXa9,b22&(fBGg;
)_=>HWCT9E2:-(^c0df,DY7V-g6.-g#GC9Ba?Q;E(JQ2&^McKH3;D)B/IUQK,^U(
4CPZB2\]C=[\P6_DV.74#=34LL-V6Hb8KD1Q90]=d=5L)LEIV>321cNUKIP/G[Ba
K??D]f/@Z.SDS@T3YcLKVV:9?G#3bSc+/^QH[eG9EAaGVHPG<88Yf=DN4/Aeae35
YKc0)=2M^4?6B1R&N5cBYZS:+IU@9Od],Q?Nd[EN3>U.>K:D#c(LQ1_#SZ:J_P2R
/a,R]Y\E:XO=-E/R;M:.a8.Fa_F=NS6^NJ=.[91B3M#YTXLQa2++MZ[)+fF36bcM
+.^<)X\/Z_-P670=Sc@YB-P]9=3ZN[\\E9(+7eD@TJc+WI+TCVdf?aQ,)2aND&;N
X^Ug7L,MW08:7SE^;3W3@gaFaC?#NDJ8[C\Naf(+)F@WHUG5L&d&dA9K#T?OB:=a
^.7XHd7C7,POGJY_(Xb([D,#PCRZ(W>8EJLafJYBTN0/XY)4=;eY9#(EI=JTb.^/
XCdZ^X(US,(SgQ>JebO:79/>[@=+aUW)>.Dc#]G]^8R@5E^&4@/<PGSX]Yc\D>dG
2N/Z>2I^+2H>4@b;9PE15+@81g^G1eT^R>&U#Z@?f/<c(:>RYU9N1@.ca92K07N&
?b8<A^S42X&147D[(IU-T-:.@9DWX34[eV+2#c,\(M=gZ4I,Ef,Cag<aJ8EeFJ9Z
&G:SN0EfX4GO,TaX9ON9MQ&C<aD=SH&\<9@54\[DM-f#+\?,(EPAKO<WHH\;1X9+
S<1#[JTC0B_#Ee7WO-76-fIN.H+YAB<<1NV+Le0B.eE5.A,H?F]6<4ER=?WS)6JP
Gd6:BZD.VEHX.GgO<XbebgMLdSS3eEO-_Y(aY\;Qg<W@gG\[I0ZR];UZ:eZgD]]H
@/IG6C,;V]WA8NAG=UC#bQ^QL?bRQ^ZD/79NNNVY=;S+?5[2(eYF)(/7CdOgP&^&
HWP;E]O.3>\?HVScaG8g@G8]I>4::H05M89.<eBX?M-VZ4]M(d[.#6G98:CY]/EP
T:#QaD?9([_\:4K#D>ccBd2QHJN1/]<=N>:>T;PSQ9Cd/Z:4Jc),;K66#gc<?W6D
RT1O.Q1/K]K&bK&+E@=Nc3CKDDRaQVB7eM4f:b0\]5/APDIYE04/b+aT)<g/)]_F
W+P?gg8-\NN-8V@4^13:Q203\-<[#EFC>5DTY_PcB-RN@2g,ZcF38V?c83aCYZ_3
RaJL6+_[MYP=V9+Q4#YW\Cg3dD1Y]C)V;/78UV8#Q<MK;X?TOTQ3ScD[(6P]6&Qg
_9D7QV0]].AS/R8bg9<27c5W8Ta#gKZ+@RaDI)(^W4#SJO8YeR[eU;fOHDD1LU3#
YNaf/IEKP5dBA#_V(8J@UH7D56fU@_6.@;0?TOTCeeO\cDcYMF&dRM+0,W;M),=.
EB\TT/)3ROe.:U_Z4+,E?GdMIH0fC)369)[8PT)XT?/dDLA74Hb9/+:K:FC^7aD_
)eM]c([MOPP6\/a0RY\c@35M^I^,S=8e;ed;U[NaQaBWT.L_=@MXS<ZW&UI:;Y6_
d;Z:a22T.H9@:B502fQX_SHH:7(#RRD6,_I6a4b]Z#+<I(H8f/#J1G<F:+W/12&e
RK.-b\:U0@dL==V-f+O-SN1LU&72:D]\AH253Bg6^205-VNJ(\8gd\UOYV=/Y^cS
5=:e\D8(b3.=[\YR&:F:X_bJ@(N<-Yd?\/XJ+Ea6/E1\Y=_JGcTAY]=aR2f9+WUg
SFcEG5=/\4-9e,1ISX[\V9ZY\[ATI6Zg&7dKUeW^e,W5J/Y=g3_K/<AI<B/geN3O
:-D9\RO+8,4,aZ?2MR7P@f@>XP+G29@<TJ:RJ;+28aAJ?Xb;JJTBV>Z+YA-C3?G,
2,;O_HZ-V;A@ZL<_FTV)/Q51)d1<?@6H9,1XcQ?=Z[\PH?#NR1CIWcT#:H5:8G];
Ne#2<&T:JQBODO+CPe-72W\c,:G8fF<1CQ37./HH&5TZ=1QNcV>+a5K7@?FSBRe;
()>ZCRK\VSS&:X35&g8YY=283b#A3O8A<S@bX42PZPV#b@:ETZIO5@I^S_QY,L6U
AUcR@_4_gQSg2_]A+#a?f.=_Q8.f\[MT<$
`endprotected
endmodule