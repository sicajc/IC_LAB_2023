`include "Usertype_FD.sv"

program automatic PATTERN_bridge(input clk, INF.PATTERN_bridge inf);
import usertype::*;

parameter DRAM_p_r = "../00_TESTBED/DRAM/dram.dat";
logic [7:0] golden_DRAM [65536+256*8-1 : 65536];
logic [16:0] addr;
logic [63:0] golden_ans;
integer patnumber = 100000;
integer i_pat, latency, total_latency, t;
// integer test1, test2, test3, test4, test5, test6, test7, test8;
initial $readmemh(DRAM_p_r, golden_DRAM);

initial begin
  reset_task;

  for (i_pat = 0; i_pat < patnumber; i_pat = i_pat+1)
    begin
        input_task;
        wait_out_valid_task;
        check_ans_task;
        $display("\033[0;34mPASS PATTERN NO.%4d,\033[m \033[0;32mexecution cycle : %3d\033[m",i_pat ,latency);
    end
  #15;
  YOU_PASS_task;
  no_out_valid_task;
end

task reset_task; begin
    inf.rst_n = 'b1;
    inf.C_in_valid = 'b0;
    inf.C_addr = 'b0;
    inf.C_data_w = 'b0;
    inf.C_r_wb = 'b0;

    total_latency = 0;

    #5; inf.rst_n = 0;
    #15; inf.rst_n = 1;

    if(inf.C_data_r !== 0) begin //out!==0
        OUO_task;
        $display ("--------------------------------------------------------------------");
        $display ("              C_data_r should be set zero after reset.              ");
        $display ("--------------------------------------------------------------------");
        repeat(5) #8;
        $finish;
    end
    if(inf.C_out_valid !== 0) begin //out!==0
        OUO_task;
        $display ("--------------------------------------------------------------------");
        $display ("             C_out_valid should be set zero after reset.            ");
        $display ("--------------------------------------------------------------------");
        repeat(5) #8;
        $finish;
    end
    if(inf.AR_VALID !== 0) begin //out!==0
        OUO_task;
        $display ("--------------------------------------------------------------------");
        $display ("             AR_VALID should be set zero after reset.               ");
        $display ("--------------------------------------------------------------------");
        repeat(5) #8;
        $finish;
    end
    if(inf.AR_ADDR !== 0) begin //out!==0
        OUO_task;
        $display ("--------------------------------------------------------------------");
        $display ("             AR_ADDR should be set zero after reset.                ");
        $display ("--------------------------------------------------------------------");
        repeat(5) #8;
        $finish;
    end
    if(inf.R_READY !== 0) begin //out!==0
        OUO_task;
        $display ("--------------------------------------------------------------------");
        $display ("             R_READY should be set zero after reset.                ");
        $display ("--------------------------------------------------------------------");
        repeat(5) #8;
        $finish;
    end
    if(inf.AW_VALID !== 0) begin //out!==0
        OUO_task;
        $display ("--------------------------------------------------------------------");
        $display ("            AW_VALID should be set zero after reset.                ");
        $display ("--------------------------------------------------------------------");
        repeat(5) #8;
        $finish;
    end
    if(inf.AW_ADDR !== 0) begin //out!==0
        OUO_task;
        $display ("--------------------------------------------------------------------");
        $display ("            AW_ADDR should be set zero after reset.                 ");
        $display ("--------------------------------------------------------------------");
        repeat(5) #8;
        $finish;
    end
    if(inf.W_VALID !== 0) begin //out!==0
        OUO_task;
        $display ("--------------------------------------------------------------------");
        $display ("            W_VALID should be set zero after reset.                 ");
        $display ("--------------------------------------------------------------------");
        repeat(5) #8;
        $finish;
    end
    if(inf.W_DATA !== 0) begin //out!==0
        OUO_task;
        $display ("--------------------------------------------------------------------");
        $display ("             W_DATA should be set zero after reset.                 ");
        $display ("--------------------------------------------------------------------");
        repeat(5) #8;
        $finish;
    end
    if(inf.B_READY !== 0) begin //out!==0
        OUO_task;
        $display ("--------------------------------------------------------------------");
        $display ("             B_READY should be set zero after reset.                ");
        $display ("--------------------------------------------------------------------");
        repeat(5) #8;
        $finish;
    end
end endtask

task input_task; begin
    t = $urandom_range(2, 10);
    repeat(1) @(negedge clk);

	// wait_out_valid_task;

    inf.C_in_valid = 'b1;
    inf.C_addr = $urandom()%255;
    inf.C_data_w[31:0] = $urandom();
    inf.C_data_w[63:32] = $urandom();
    inf.C_r_wb = $urandom()%2;

    @(negedge clk);

    inf.C_in_valid = 'b0;
    addr = 17'h10000+inf.C_addr*8;

    if (inf.C_r_wb==0) begin
    	golden_DRAM[addr+7] = inf.C_data_w[63:56];
    	golden_DRAM[addr+6] = inf.C_data_w[55:48];
    	golden_DRAM[addr+5] = inf.C_data_w[47:40];
    	golden_DRAM[addr+4] = inf.C_data_w[39:32];
    	golden_DRAM[addr+3] = inf.C_data_w[31:24];
    	golden_DRAM[addr+2] = inf.C_data_w[23:16];
    	golden_DRAM[addr+1] = inf.C_data_w[15:8];
    	golden_DRAM[addr] = inf.C_data_w[7:0];
    end

    golden_ans = {golden_DRAM[addr+7],
    			  golden_DRAM[addr+6],
    			  golden_DRAM[addr+5],
    			  golden_DRAM[addr+4],
    			  golden_DRAM[addr+3],
    			  golden_DRAM[addr+2],
    			  golden_DRAM[addr+1],
    			  golden_DRAM[addr]};

end endtask

task wait_out_valid_task; begin
    latency = 0;
    while(inf.C_out_valid !== 1'b1) begin
        latency = latency + 1;

        if( latency == 1000) begin
        	OUO_task;
            $display ("--------------------------------------------------------------------");
            $display ("         The execution latency is limited in 1000 cycles.           ");
            $display ("--------------------------------------------------------------------");
            repeat(5) #8;
            $finish;
        end
        @(negedge clk);
    end
    total_latency = total_latency + latency;
end endtask

task no_out_valid_task; begin
    latency = 0;
    while(inf.C_out_valid === 1'b0) begin
        latency = latency + 1;

        if( latency == 1000) begin
            $finish;
        end
        @(negedge clk);
    end
    OUO_task;
    $display ("--------------------------------------------------------------------------");
    $display ("The out_valid should set to low even if you pass all of the TA’s patterns.");
    $display ("--------------------------------------------------------------------------");
    $finish;
end endtask

task check_ans_task; begin
	if (inf.C_r_wb) begin
    	if (inf.C_data_r!==golden_ans) begin
    	    show_ans_task;
    	    repeat(5) #8;
    	    $finish;
    	end
	end
end endtask

task show_ans_task; begin
    OUO_task;
    $display ("ADDRESS: %d",inf.C_addr);
    $display ("YOUR   : %2h %2h %2h %2h_%2h %2h %2h %2h",inf.C_data_r[63:56]
                                                        ,inf.C_data_r[55:48]
                                                        ,inf.C_data_r[47:40]
                                                        ,inf.C_data_r[39:32]
                                                        ,inf.C_data_r[31:24]
                                                        ,inf.C_data_r[23:16]
                                                        ,inf.C_data_r[15:8]
                                                        ,inf.C_data_r[7:0]);
    $display ("GOLDEN : %2h %2h %2h %2h_%2h %2h %2h %2h",golden_ans[63:56]
                                                        ,golden_ans[55:48]
                                                        ,golden_ans[47:40]
                                                        ,golden_ans[39:32]
                                                        ,golden_ans[31:24]
                                                        ,golden_ans[23:16]
                                                        ,golden_ans[15:8]
                                                        ,golden_ans[7:0]);

end endtask

task OUO_task; begin
  $display ("\033[49m  \033[38;2;186;167;118;49m \033[38;2;53;38;21;48;2;52;30;18m \033[38;2;16;15;8;48;2;20;15;14m \033[38;2;19;19;22;48;2;19;18;19m \033[38;2;13;13;18;48;2;17;16;17m \033[38;2;11;11;16;48;2;14;13;14m \033[38;2;13;13;20;48;2;16;15;17m \033[38;2;11;10;18;48;2;14;13;16m \033[38;2;13;12;15;48;2;14;12;15m \033[38;2;14;12;13;48;2;14;13;14m \033[38;2;12;11;11;48;2;13;11;11m \033[38;2;16;15;15;48;2;16;15;16m \033[38;2;14;10;17;48;2;13;9;15m \033[38;2;14;10;17;48;2;12;8;16m \033[38;2;10;10;15;48;2;11;11;17m \033[38;2;3;9;14;48;2;7;8;15m \033[38;2;6;7;13;48;2;8;11;16m \033[38;2;9;10;16;48;2;12;11;17m \033[38;2;9;10;16;48;2;9;9;15m \033[38;2;10;10;15;48;2;10;10;16m \033[38;2;10;11;17;48;2;11;13;18m \033[38;2;4;8;17;48;2;4;9;17m \033[48;2;3;7;17m \033[38;2;3;7;17;48;2;3;8;17m \033[38;2;3;7;17;48;2;6;10;19m \033[38;2;3;7;17;48;2;6;10;20m \033[38;2;2;6;16;48;2;2;6;15m \033[38;2;4;10;15;48;2;5;11;15m \033[38;2;6;13;17;48;2;9;13;17m \033[38;2;4;9;13;48;2;9;9;14m \033[38;2;13;11;16;48;2;13;12;17m \033[38;2;20;18;26;48;2;21;17;25m \033[38;2;21;18;26;48;2;19;16;23m \033[38;2;20;18;25;48;2;18;17;23m \033[38;2;18;16;22;48;2;15;12;18m \033[38;2;15;12;17;48;2;12;9;15m \033[38;2;16;14;19;48;2;18;16;21m \033[38;2;18;16;22;48;2;19;16;22m \033[m");
  $display ("\033[49m \033[38;2;138;86;52;49m \033[38;2;117;74;55;48;2;137;96;58m \033[38;2;35;23;15;48;2;39;26;11m \033[38;2;16;17;12;48;2;15;17;8m \033[38;2;19;20;19;48;2;19;19;22m \033[38;2;13;14;17;48;2;13;13;18m \033[38;2;9;8;13;48;2;10;10;18m \033[38;2;9;8;15;48;2;12;13;20m \033[38;2;9;8;15;48;2;10;9;16m \033[38;2;13;11;14;48;2;14;10;15m \033[48;2;15;14;14m \033[38;2;12;11;11;48;2;12;10;11m \033[38;2;15;13;14;48;2;15;13;13m \033[38;2;16;13;19;48;2;16;12;18m \033[38;2;17;13;20;48;2;16;11;18m \033[38;2;10;8;14;48;2;9;8;14m \033[38;2;1;6;11;48;2;1;7;12m \033[38;2;4;7;12;48;2;2;6;11m \033[38;2;4;8;13;48;2;3;9;14m \033[38;2;0;5;9;48;2;5;10;14m \033[38;2;5;7;11;48;2;8;10;16m \033[38;2;9;9;14;48;2;10;10;17m \033[38;2;6;8;15;48;2;4;8;16m \033[38;2;5;7;15;48;2;3;7;17m \033[38;2;4;6;14;48;2;3;7;17m \033[38;2;6;6;15;48;2;3;7;17m \033[38;2;7;8;16;48;2;3;7;17m \033[38;2;4;5;12;48;2;1;5;15m \033[38;2;6;6;17;48;2;3;9;14m \033[38;2;8;7;17;48;2;7;12;17m \033[38;2;6;6;16;48;2;5;8;13m \033[38;2;7;8;16;48;2;9;7;13m \033[38;2;17;17;20;48;2;20;18;25m \033[38;2;24;22;27;48;2;23;19;27m \033[38;2;21;18;25;48;2;22;19;26m \033[38;2;17;14;20;48;2;18;15;21m \033[38;2;13;9;15;48;2;15;12;19m \033[38;2;14;11;16;48;2;16;13;19m \033[38;2;12;13;18;48;2;18;16;22m \033[m");
  $display ("\033[49m \033[38;2;124;66;44;48;2;123;71;42m \033[38;2;115;77;76;48;2;111;72;63m \033[38;2;27;21;14;48;2;32;22;13m \033[38;2;22;19;16;48;2;18;16;10m \033[38;2;22;26;17;48;2;18;23;15m \033[38;2;19;17;14;48;2;13;16;12m \033[38;2;8;7;12;48;2;7;7;13m \033[38;2;8;7;13;48;2;8;8;12m \033[38;2;9;9;13;48;2;9;9;14m \033[38;2;12;9;13;48;2;13;11;13m \033[38;2;14;12;12;48;2;14;13;13m \033[48;2;14;12;13m \033[38;2;17;14;18;48;2;17;13;17m \033[38;2;21;17;24;48;2;20;16;23m \033[38;2;22;18;26;48;2;21;17;25m \033[38;2;15;10;18;48;2;13;9;15m \033[38;2;4;6;11;48;2;2;5;10m \033[38;2;8;7;13;48;2;7;7;13m \033[38;2;7;9;14;48;2;6;8;13m \033[38;2;1;6;10;48;2;1;5;9m \033[38;2;5;6;10;48;2;4;5;9m \033[38;2;8;8;13;48;2;8;7;11m \033[38;2;10;10;15;48;2;9;8;13m \033[38;2;9;8;15;48;2;7;7;13m \033[38;2;7;7;13;48;2;5;4;10m \033[38;2;9;8;15;48;2;7;6;13m \033[38;2;14;14;20;48;2;11;11;17m \033[38;2;12;11;18;48;2;8;7;14m \033[38;2;10;8;18;48;2;9;7;18m \033[38;2;9;7;18;48;2;9;6;18m \033[48;2;7;6;17m \033[38;2;8;10;18;48;2;8;11;19m \033[38;2;13;12;16;48;2;13;13;17m \033[38;2;21;19;23;48;2;22;20;25m \033[38;2;24;21;28;48;2;22;20;27m \033[38;2;13;10;17;48;2;15;12;18m \033[38;2;13;10;18;48;2;13;10;16m \033[38;2;9;7;14;48;2;12;8;16m \033[38;2;9;9;15;48;2;10;10;17m \033[m");
  $display ("\033[38;2;123;66;19;48;2;137;78;20m \033[38;2;130;80;56;48;2;129;69;54m \033[38;2;78;44;57;48;2;101;59;58m \033[38;2;47;32;29;48;2;25;16;14m \033[38;2;84;69;68;48;2;45;37;38m \033[38;2;85;70;72;48;2;45;41;36m \033[38;2;64;51;44;48;2;30;25;23m \033[38;2;31;29;29;48;2;16;13;20m \033[38;2;13;14;13;48;2;9;9;15m \033[38;2;11;7;12;48;2;9;9;13m \033[38;2;12;8;13;48;2;10;6;11m \033[38;2;14;12;13;48;2;14;12;12m \033[38;2;14;12;12;48;2;15;14;13m \033[38;2;16;12;15;48;2;18;16;19m \033[38;2;20;15;19;48;2;22;18;22m \033[38;2;21;17;19;48;2;22;18;24m \033[38;2;18;14;20;48;2;17;13;20m \033[38;2;14;14;20;48;2;11;12;18m \033[38;2;14;12;18;48;2;10;9;16m \033[38;2;12;10;17;48;2;8;8;12m \033[38;2;10;9;15;48;2;2;7;10m \033[38;2;9;8;14;48;2;5;7;13m \033[38;2;15;14;20;48;2;10;10;16m \033[38;2;19;16;23;48;2;12;11;18m \033[38;2;15;11;19;48;2;10;9;15m \033[38;2;13;9;16;48;2;9;8;13m \033[38;2;14;10;17;48;2;11;9;15m \033[38;2;24;22;30;48;2;16;15;22m \033[38;2;21;18;26;48;2;16;15;22m \033[38;2;12;8;20;48;2;11;9;20m \033[38;2;9;6;19;48;2;9;6;18m \033[38;2;7;5;17;48;2;7;5;16m \033[38;2;13;12;18;48;2;11;12;18m \033[38;2;18;14;21;48;2;16;13;18m \033[38;2;26;19;24;48;2;23;18;24m \033[38;2;33;27;35;48;2;29;24;32m \033[38;2;12;12;25;48;2;14;13;21m \033[38;2;8;7;19;48;2;10;9;16m \033[38;2;6;6;18;48;2;8;8;16m \033[38;2;3;6;17;48;2;6;8;15m \033[m");
  $display ("\033[38;2;133;83;44;48;2;124;76;34m \033[38;2;111;73;50;48;2;115;75;55m \033[38;2;62;37;28;48;2;43;23;22m \033[38;2;99;85;67;48;2;73;62;49m \033[38;2;111;93;73;48;2;104;91;76m \033[38;2;110;90;74;48;2;108;89;78m \033[38;2;102;81;68;48;2;98;83;66m \033[38;2;94;74;64;48;2;80;73;64m \033[38;2;76;60;56;48;2;46;38;36m \033[38;2;61;44;46;48;2;28;19;19m \033[38;2;50;36;35;48;2;25;19;21m \033[38;2;47;32;35;48;2;25;20;22m \033[38;2;46;35;35;48;2;23;17;19m \033[38;2;42;32;35;48;2;19;14;15m \033[38;2;29;21;27;48;2;17;13;16m \033[38;2;18;13;16;48;2;19;12;16m \033[38;2;21;17;21;48;2;20;14;21m \033[38;2;20;18;21;48;2;16;15;19m \033[38;2;20;16;21;48;2;17;14;19m \033[38;2;21;15;24;48;2;18;14;19m \033[38;2;20;15;22;48;2;14;10;18m \033[38;2;16;11;18;48;2;13;9;17m \033[38;2;15;11;17;48;2;15;12;19m \033[48;2;18;15;21m \033[38;2;20;16;23;48;2;18;16;22m \033[38;2;21;16;22;48;2;18;14;20m \033[38;2;24;16;24;48;2;19;15;22m \033[38;2;45;40;53;48;2;31;28;40m \033[38;2;27;21;33;48;2;25;21;33m \033[38;2;14;10;22;48;2;13;9;20m \033[38;2;9;9;20;48;2;8;7;20m \033[38;2;8;9;19;48;2;8;7;18m \033[38;2;14;11;23;48;2;14;12;23m \033[38;2;17;12;23;48;2;18;15;23m \033[38;2;27;22;30;48;2;28;23;30m \033[38;2;26;22;29;48;2;32;26;35m \033[38;2;10;9;20;48;2;13;11;22m \033[38;2;4;6;19;48;2;7;6;19m \033[38;2;3;6;17;48;2;5;5;18m \033[38;2;1;4;15;48;2;3;4;16m \033[m");
  $display ("\033[38;2;125;82;48;48;2;135;90;60m \033[38;2;101;60;41;48;2;107;70;52m \033[38;2;108;80;67;48;2;83;61;51m \033[38;2;114;95;72;48;2;112;94;76m \033[38;2;108;86;64;48;2;111;90;74m \033[38;2;96;69;50;48;2;99;75;61m \033[38;2;81;51;37;48;2;91;65;53m \033[38;2;65;43;29;48;2;83;61;48m \033[38;2;46;30;19;48;2;67;51;43m \033[38;2;34;17;14;48;2;64;47;49m \033[38;2;37;23;21;48;2;60;46;47m \033[38;2;38;28;29;48;2;58;42;41m \033[38;2;57;44;48;48;2;60;43;43m \033[38;2;70;51;57;48;2;64;48;49m \033[38;2;77;58;61;48;2;59;45;44m \033[38;2;86;62;66;48;2;48;36;32m \033[38;2;96;71;73;48;2;50;37;36m \033[38;2;103;72;71;48;2;42;26;27m \033[38;2;107;76;71;48;2;41;25;28m \033[38;2;110;80;76;48;2;47;31;38m \033[38;2;100;71;72;48;2;34;19;25m \033[38;2;71;45;43;48;2;22;11;13m \033[38;2;54;35;32;48;2;19;14;16m \033[38;2;48;35;37;48;2;21;17;22m \033[38;2;30;18;18;48;2;21;16;19m \033[38;2;36;25;29;48;2;24;15;20m \033[38;2;49;32;37;48;2;32;21;28m \033[38;2;48;34;36;48;2;46;35;47m \033[38;2;28;19;23;48;2;26;18;27m \033[38;2;19;15;22;48;2;16;11;21m \033[38;2;13;11;20;48;2;9;9;20m \033[38;2;9;10;21;48;2;8;9;18m \033[38;2;11;9;21;48;2;10;6;19m \033[38;2;16;13;22;48;2;14;8;18m \033[38;2;21;17;26;48;2;21;16;24m \033[38;2;14;11;18;48;2;19;17;23m \033[38;2;8;7;16;48;2;8;8;18m \033[38;2;6;6;18;48;2;4;7;18m \033[38;2;5;7;16;48;2;2;6;17m \033[38;2;3;8;14;48;2;1;6;14m \033[m");
  $display ("\033[38;2;119;78;48;48;2;129;86;51m \033[38;2;114;74;55;48;2;103;60;42m \033[38;2;125;99;77;48;2;122;94;78m \033[38;2;116;94;67;48;2;115;93;68m \033[38;2;109;88;53;48;2;106;89;55m \033[38;2;105;82;53;48;2;98;78;51m \033[38;2;98;74;51;48;2;81;58;37m \033[38;2;81;61;45;48;2;57;39;22m \033[38;2;67;50;38;48;2;39;21;11m \033[38;2;57;39;35;48;2;32;16;10m \033[38;2;39;30;30;48;2;13;6;6m \033[38;2;12;7;6;48;2;0;1;0m \033[38;2;12;13;11;48;2;19;21;28m \033[38;2;92;92;97;48;2;78;72;83m \033[38;2;97;95;99;48;2;74;58;61m \033[38;2;68;55;53;48;2;85;62;66m \033[38;2;99;67;67;48;2;101;72;73m \033[38;2;119;79;74;48;2;122;86;81m \033[38;2;123;85;74;48;2;125;90;80m \033[38;2;127;88;73;48;2;132;93;88m \033[38;2;144;102;90;48;2;140;98;98m \033[38;2;155;109;99;48;2;136;95;92m \033[38;2;162;118;108;48;2;130;93;85m \033[38;2;162;121;110;48;2;111;75;68m \033[38;2;163;121;112;48;2;85;44;35m \033[38;2;157;112;103;48;2;93;55;49m \033[38;2;147;105;103;48;2;95;65;60m \033[38;2;118;87;86;48;2;67;51;49m \033[38;2;96;68;68;48;2;44;29;27m \033[38;2;81;60;60;48;2;37;24;28m \033[38;2;64;45;42;48;2;25;15;22m \033[38;2;68;49;47;48;2;19;13;20m \033[38;2;69;51;51;48;2;28;21;28m \033[38;2;64;48;52;48;2;26;20;29m \033[38;2;51;42;48;48;2;29;23;33m \033[38;2;26;15;23;48;2;20;14;22m \033[38;2;20;13;19;48;2;12;7;14m \033[38;2;19;15;21;48;2;9;7;11m \033[38;2;20;15;22;48;2;12;9;16m \033[38;2;16;13;20;48;2;11;11;18m \033[m");
  $display ("\033[38;2;125;89;47;48;2;121;84;47m \033[38;2;130;96;66;48;2;122;89;66m \033[38;2;135;106;77;48;2;127;102;71m \033[38;2;131;100;68;48;2;123;94;68m \033[38;2;129;93;64;48;2;123;88;59m \033[38;2;124;85;58;48;2;118;84;56m \033[38;2;118;83;59;48;2;109;79;57m \033[38;2;111;79;61;48;2;98;72;56m \033[38;2;104;71;61;48;2;89;65;50m \033[38;2;93;65;56;48;2;79;54;43m \033[38;2;85;63;55;48;2;64;46;39m \033[38;2;81;59;52;48;2;51;37;31m \033[38;2;79;57;49;48;2;50;38;30m \033[38;2;72;51;43;48;2;59;45;40m \033[38;2;72;49;43;48;2;55;38;37m \033[38;2;83;55;52;48;2;54;30;27m \033[38;2;99;67;62;48;2;92;60;59m \033[38;2;105;70;61;48;2;113;76;72m \033[38;2;107;72;53;48;2;114;78;66m \033[38;2;119;82;61;48;2;118;84;64m \033[38;2;145;99;83;48;2;147;101;87m \033[38;2;157;111;98;48;2;158;113;101m \033[38;2;172;128;117;48;2;173;129;123m \033[38;2;173;130;124;48;2;173;131;124m \033[38;2;173;133;124;48;2;171;130;123m \033[38;2;161;118;105;48;2;165;123;112m \033[38;2;144;103;95;48;2;151;108;101m \033[38;2;104;78;70;48;2;122;87;84m \033[38;2;44;29;25;48;2;102;75;70m \033[38;2;30;13;19;48;2;84;62;56m \033[38;2;53;37;46;48;2;80;58;48m \033[38;2;78;63;65;48;2;84;63;57m \033[38;2;80;63;59;48;2;88;64;61m \033[38;2;77;60;57;48;2;82;63;62m \033[38;2;76;58;56;48;2;68;51;52m \033[38;2;77;61;63;48;2;41;27;31m \033[38;2;88;63;64;48;2;42;28;31m \033[38;2;100;70;67;48;2;52;35;36m \033[38;2;109;78;70;48;2;55;34;41m \033[38;2;109;74;63;48;2;37;16;19m \033[m");
  $display ("\033[38;2;140;120;80;48;2;130;91;52m \033[38;2;145;118;85;48;2;144;108;72m \033[38;2;154;121;89;48;2;150;119;85m \033[38;2;154;119;86;48;2;149;115;81m \033[38;2;158;118;85;48;2;149;111;79m \033[38;2;162;120;92;48;2;144;102;75m \033[38;2;161;120;90;48;2;135;96;70m \033[38;2;161;119;93;48;2;129;88;71m \033[38;2;161;117;92;48;2;119;80;65m \033[38;2;148;102;75;48;2;113;75;60m \033[38;2;130;81;61;48;2;109;70;59m \033[38;2;121;73;59;48;2;105;66;59m \033[38;2;116;73;58;48;2;98;61;55m \033[38;2;115;73;60;48;2;94;63;53m \033[38;2;112;77;64;48;2;95;66;56m \033[38;2;111;77;65;48;2;99;70;58m \033[38;2;110;77;62;48;2;102;70;60m \033[38;2;111;79;57;48;2;105;72;57m \033[38;2;135;97;68;48;2;112;76;53m \033[38;2;184;145;121;48;2;129;91;65m \033[38;2;219;188;177;48;2;155;110;90m \033[38;2;219;188;178;48;2;165;119;101m \033[38;2;184;140;117;48;2;170;126;107m \033[38;2;174;125;106;48;2;170;125;112m \033[38;2;167;124;114;48;2;166;124;115m \033[38;2;154;109;98;48;2;154;112;99m \033[38;2;144;103;93;48;2;143;104;96m \033[38;2;123;85;83;48;2;68;49;38m \033[38;2;67;47;46;48;2;5;1;1m \033[38;2;35;23;30;48;2;3;0;7m \033[38;2;42;33;41;48;2;31;27;38m \033[38;2;106;91;102;48;2;104;98;107m \033[38;2;114;92;97;48;2;105;93;92m \033[38;2;86;63;64;48;2;78;61;59m \033[38;2;62;40;39;48;2;62;42;40m \033[38;2;61;39;36;48;2;61;41;40m \033[38;2;91;57;52;48;2;84;58;53m \033[38;2;112;69;60;48;2;104;68;60m \033[38;2;119;73;57;48;2;113;75;61m \033[38;2;127;77;57;48;2;124;84;66m \033[m");
  $display ("\033[38;2;145;117;80;48;2;147;119;84m \033[38;2;142;111;78;48;2;144;113;80m \033[38;2;147;113;80;48;2;148;114;80m \033[38;2;154;116;83;48;2;153;115;82m \033[38;2;165;120;91;48;2;161;118;88m \033[38;2;177;128;102;48;2;169;123;96m \033[38;2;184;136;114;48;2;172;128;101m \033[38;2;190;144;121;48;2;175;131;107m \033[38;2;192;147;122;48;2;179;136;113m \033[38;2;192;148;121;48;2;173;129;103m \033[38;2;189;144;120;48;2;159;109;86m \033[38;2;172;121;101;48;2;146;95;78m \033[38;2;154;102;79;48;2;140;90;74m \033[38;2;150;101;77;48;2;136;92;73m \033[38;2;145;99;73;48;2;134;92;71m \033[38;2;143;98;68;48;2;130;90;67m \033[38;2;155;110;78;48;2;130;91;66m \033[38;2;183;138;109;48;2;143;97;71m \033[38;2;205;167;134;48;2;180;138;109m \033[38;2;231;205;181;48;2;216;189;168m \033[38;2;252;247;243;48;2;242;233;229m \033[38;2;247;234;227;48;2;240;225;219m \033[38;2;238;214;200;48;2;221;186;167m \033[38;2;221;180;161;48;2;190;136;115m \033[38;2;194;142;126;48;2;178;127;116m \033[38;2;181;129;111;48;2;167;118;106m \033[38;2;166;119;105;48;2;151;104;95m \033[38;2;149;102;97;48;2;132;87;86m \033[38;2;130;85;82;48;2;111;71;69m \033[38;2;123;81;82;48;2;102;68;72m \033[38;2;126;86;79;48;2;99;68;68m \033[38;2;131;92;82;48;2;101;71;65m \033[38;2;138;100;87;48;2;107;77;72m \033[38;2;147;110;93;48;2;116;83;73m \033[38;2;155;115;91;48;2;121;86;70m \033[38;2;162;119;96;48;2;125;88;71m \033[38;2;164;121;98;48;2;133;92;77m \033[38;2;168;120;99;48;2;143;97;85m \033[38;2;171;120;95;48;2;146;98;79m \033[38;2;175;123;95;48;2;153;102;80m \033[m");
  $display ("\033[38;2;138;106;81;48;2;140;110;79m \033[38;2;140;106;81;48;2;141;109;80m \033[38;2;149;111;84;48;2;149;112;82m \033[38;2;161;119;94;48;2;158;117;90m \033[38;2;170;125;100;48;2;168;122;96m \033[38;2;179;129;102;48;2;178;128;100m \033[38;2;186;137;110;48;2;187;136;111m \033[38;2;196;145;119;48;2;194;145;121m \033[38;2;202;154;126;48;2;198;152;124m \033[38;2;206;160;131;48;2;202;156;127m \033[38;2;206;162;132;48;2;201;157;131m \033[38;2;204;162;134;48;2;196;151;126m \033[38;2;197;154;129;48;2;180;132;107m \033[38;2;175;126;99;48;2;165;118;93m \033[38;2;158;106;78;48;2;155;108;82m \033[38;2;161;115;78;48;2;154;110;76m \033[38;2;184;141;103;48;2;177;132;98m \033[38;2;218;179;148;48;2;199;156;123m \033[38;2;237;208;184;48;2;220;186;156m \033[38;2;246;232;215;48;2;242;224;203m \033[38;2;254;251;249;48;2;253;252;250m \033[38;2;250;239;229;48;2;249;238;228m \033[38;2;245;228;213;48;2;243;224;214m \033[38;2;240;217;202;48;2;237;212;197m \033[38;2;229;194;178;48;2;214;169;148m \033[38;2;209;160;138;48;2;195;143;121m \033[38;2;199;152;135;48;2;186;138;121m \033[38;2;183;132;120;48;2;168;119;111m \033[38;2;175;124;110;48;2;153;104;95m \033[38;2;164;116;99;48;2;142;96;87m \033[38;2;161;113;95;48;2;145;100;87m \033[38;2;164;117;99;48;2;151;105;90m \033[38;2;170;124;107;48;2;157;114;97m \033[38;2;182;138;118;48;2;168;128;107m \033[38;2;190;145;120;48;2;174;133;105m \033[38;2;197;150;122;48;2;181;136;107m \033[38;2;203;158;128;48;2;186;140;110m \033[38;2;213;176;148;48;2;192;146;117m \033[38;2;219;185;158;48;2;200;160;130m \033[38;2;218;184;156;48;2;200;158;124m \033[m");
  $display ("\033[38;2;136;109;85;48;2;134;103;81m \033[38;2;140;110;86;48;2;138;106;82m \033[38;2;150;115;87;48;2;149;112;84m \033[38;2;162;123;96;48;2;162;122;98m \033[38;2;172;131;108;48;2;173;129;106m \033[38;2;183;139;118;48;2;183;136;113m \033[38;2;193;148;125;48;2;192;145;121m \033[38;2;199;152;126;48;2;199;150;125m \033[38;2;205;157;128;48;2;204;156;128m \033[38;2;210;165;135;48;2;208;163;133m \033[38;2;211;168;138;48;2;208;165;135m \033[38;2;208;168;138;48;2;207;166;137m \033[38;2;200;159;133;48;2;201;159;135m \033[38;2;168;112;79;48;2;175;119;89m \033[38;2;173;126;95;48;2;153;93;60m \033[38;2;197;170;143;48;2;173;131;96m \033[38;2;222;197;171;48;2;212;178;146m \033[38;2;238;213;195;48;2;236;205;180m \033[38;2;242;223;204;48;2;245;224;208m \033[38;2;248;238;227;48;2;252;247;240m \033[38;2;253;249;246;48;2;254;251;249m \033[38;2;252;242;237;48;2;250;240;230m \033[38;2;248;232;221;48;2;246;229;215m \033[38;2;242;215;198;48;2;238;212;195m \033[38;2;234;202;184;48;2;234;203;185m \033[38;2;219;171;143;48;2;217;172;150m \033[38;2;207;160;135;48;2;205;160;138m \033[38;2;197;146;122;48;2;190;137;120m \033[38;2;193;142;118;48;2;186;133;115m \033[38;2;195;144;121;48;2;183;130;111m \033[38;2;198;150;128;48;2;181;126;108m \033[38;2;197;149;127;48;2;182;127;109m \033[38;2;201;155;133;48;2;188;134;117m \033[38;2;210;168;148;48;2;200;152;132m \033[38;2;219;176;151;48;2;210;164;141m \033[38;2;222;179;150;48;2;214;169;140m \033[38;2;227;187;155;48;2;220;180;150m \033[38;2;230;194;163;48;2;226;192;163m \033[38;2;232;200;173;48;2;228;195;168m \033[38;2;232;202;175;48;2;227;194;167m \033[m");
  $display ("\033[38;2;138;113;90;48;2;137;113;89m \033[38;2;143;116;92;48;2;143;115;90m \033[38;2;154;121;95;48;2;153;118;91m \033[38;2;162;124;99;48;2;161;122;96m \033[38;2;169;127;105;48;2;170;128;107m \033[38;2;177;132;111;48;2;180;135;116m \033[38;2;186;139;117;48;2;190;145;123m \033[38;2;194;145;120;48;2;197;150;124m \033[38;2;203;155;127;48;2;204;156;128m \033[38;2;211;166;137;48;2;211;166;136m \033[38;2;213;170;141;48;2;213;170;140m \033[38;2;210;171;142;48;2;209;169;138m \033[38;2;194;146;115;48;2;197;151;124m \033[38;2;186;141;116;48;2;190;143;117m \033[38;2;167;117;90;48;2;191;152;126m \033[38;2;164;121;94;48;2;195;164;135m \033[38;2;192;150;123;48;2;216;188;159m \033[38;2;219;177;156;48;2;234;206;186m \033[38;2;229;194;171;48;2;239;211;192m \033[38;2;234;206;187;48;2;243;221;203m \033[38;2;239;214;196;48;2;247;231;218m \033[38;2;239;213;196;48;2;249;232;222m \033[38;2;238;211;196;48;2;247;229;216m \033[38;2;238;209;195;48;2;243;217;202m \033[38;2;238;209;195;48;2;236;206;190m \033[38;2;221;177;153;48;2;218;169;143m \033[38;2;204;151;127;48;2;205;154;129m \033[38;2;206;156;132;48;2;201;152;128m \033[38;2;215;167;143;48;2;204;156;132m \033[38;2;219;175;154;48;2;210;166;146m \033[38;2;222;179;158;48;2;212;170;150m \033[38;2;223;181;160;48;2;211;167;144m \033[38;2;226;184;165;48;2;213;170;148m \033[38;2;228;190;169;48;2;221;182;162m \033[38;2;229;190;168;48;2;225;185;162m \033[38;2;229;189;165;48;2;226;186;159m \033[38;2;227;186;159;48;2;227;187;158m \033[38;2;226;185;153;48;2;228;189;157m \033[38;2;225;185;152;48;2;229;191;159m \033[38;2;225;186;153;48;2;230;196;166m \033[m");
  $display ("\033[38;2;131;105;83;48;2;135;110;85m \033[38;2;136;106;82;48;2;140;112;88m \033[38;2;143;107;81;48;2;150;116;89m \033[38;2;152;111;84;48;2;160;120;96m \033[38;2;160;115;90;48;2;166;124;100m \033[38;2;166;118;94;48;2;173;127;105m \033[38;2;176;127;100;48;2;182;134;111m \033[38;2;188;137;111;48;2;190;140;115m \033[38;2;197;146;119;48;2;201;151;124m \033[38;2;205;157;130;48;2;208;162;135m \033[38;2;208;163;142;48;2;211;167;143m \033[38;2;202;157;141;48;2;210;170;147m \033[38;2;135;73;53;48;2;177;123;96m \033[38;2;126;76;56;48;2;155;107;81m \033[38;2;104;64;52;48;2;106;57;39m \033[38;2;86;45;36;48;2;93;54;42m \033[38;2;100;57;40;48;2;141;104;88m \033[38;2;145;95;76;48;2;180;130;114m \033[38;2;164;109;91;48;2;199;150;128m \033[38;2;166;107;90;48;2;210;168;147m \033[38;2;161;109;93;48;2;210;167;147m \033[38;2;116;72;60;48;2;213;167;148m \033[38;2;83;48;42;48;2;213;166;150m \033[38;2;165;129;116;48;2;223;183;164m \033[38;2;223;180;152;48;2;235;203;185m \033[38;2;227;191;164;48;2;229;195;177m \033[38;2;211;160;136;48;2;205;153;129m \033[38;2;216;171;150;48;2;212;165;139m \033[38;2;223;181;159;48;2;220;174;152m \033[38;2;227;187;166;48;2;224;183;162m \033[38;2;229;191;169;48;2;227;188;166m \033[38;2;230;192;169;48;2;228;190;168m \033[38;2;230;190;167;48;2;231;192;170m \033[38;2;228;188;164;48;2;230;192;170m \033[38;2;228;187;163;48;2;230;191;168m \033[38;2;225;183;158;48;2;228;188;164m \033[38;2;221;175;145;48;2;225;182;155m \033[38;2;218;171;140;48;2;222;178;146m \033[38;2;218;171;139;48;2;221;178;145m \033[38;2;217;170;138;48;2;221;177;144m \033[m");
  $display ("\033[38;2;125;100;83;48;2;128;102;83m \033[38;2;132;102;81;48;2;135;104;82m \033[38;2;139;103;79;48;2;142;105;81m \033[38;2;147;106;80;48;2;151;109;82m \033[38;2;155;111;84;48;2;157;111;85m \033[38;2;159;113;88;48;2;163;113;89m \033[38;2;164;118;93;48;2;172;119;97m \033[38;2;171;124;99;48;2;184;131;106m \033[38;2;178;131;106;48;2;192;140;112m \033[38;2;186;143;121;48;2;199;150;124m \033[38;2;190;151;129;48;2;203;159;136m \033[38;2;184;145;130;48;2;197;152;138m \033[38;2;161;110;96;48;2;135;75;60m \033[38;2;138;93;78;48;2;126;77;63m \033[38;2;132;91;83;48;2;114;76;67m \033[38;2;137;96;86;48;2;117;81;73m \033[38;2;143;101;91;48;2;124;85;67m \033[38;2;149;109;99;48;2;136;94;76m \033[38;2;147;105;94;48;2;147;102;85m \033[38;2;147;103;89;48;2;151;102;86m \033[38;2;151;105;90;48;2;142;96;83m \033[38;2;152;106;92;48;2;109;70;63m \033[38;2;152;103;94;48;2;58;27;24m \033[38;2;151;96;85;48;2;75;37;29m \033[38;2;172;114;99;48;2;185;133;110m \033[38;2;202;144;116;48;2;215;164;132m \033[38;2;220;178;154;48;2;216;169;144m \033[38;2;224;183;158;48;2;220;177;155m \033[38;2;225;184;159;48;2;224;183;159m \033[38;2;226;186;161;48;2;227;187;164m \033[38;2;228;188;164;48;2;229;191;167m \033[38;2;228;187;163;48;2;229;191;167m \033[38;2;225;183;156;48;2;227;186;160m \033[38;2;224;181;154;48;2;226;184;157m \033[38;2;224;182;156;48;2;226;184;158m \033[38;2;223;181;154;48;2;223;180;154m \033[38;2;219;174;146;48;2;219;173;144m \033[38;2;216;168;140;48;2;217;169;139m \033[38;2;213;165;136;48;2;215;167;138m \033[38;2;211;160;132;48;2;214;166;136m \033[m");
  $display ("\033[38;2;113;89;72;48;2;120;96;80m \033[38;2;123;96;80;48;2;126;98;80m \033[38;2;128;94;76;48;2;133;98;76m \033[38;2;133;95;74;48;2;139;100;76m \033[38;2;137;96;74;48;2;146;104;80m \033[38;2;141;100;77;48;2;152;110;84m \033[38;2;142;104;81;48;2;153;112;85m \033[38;2;146;109;87;48;2;156;117;90m \033[38;2;144;108;93;48;2;163;124;99m \033[38;2;138;102;89;48;2;169;130;107m \033[38;2;131;91;80;48;2;168;129;105m \033[38;2;132;90;81;48;2;164;125;107m \033[38;2;140;98;95;48;2;163;124;106m \033[38;2;140;99;93;48;2;153;115;104m \033[38;2;133;90;80;48;2;143;105;94m \033[38;2;139;93;85;48;2;146;107;96m \033[38;2;151;109;102;48;2;150;112;103m \033[38;2;155;110;106;48;2;153;114;105m \033[38;2;148;101;95;48;2;147;106;95m \033[38;2;153;106;98;48;2;146;104;90m \033[38;2;165;122;114;48;2;157;115;98m \033[38;2;176;138;127;48;2;161;118;103m \033[38;2;181;144;131;48;2;164;118;105m \033[38;2;180;141;130;48;2;169;120;111m \033[38;2;187;139;125;48;2;176;118;106m \033[38;2;217;179;157;48;2;197;140;113m \033[38;2;234;207;193;48;2;229;197;180m \033[38;2;229;195;172;48;2;226;189;163m \033[38;2;225;184;158;48;2;226;185;159m \033[38;2;224;182;157;48;2;226;185;159m \033[38;2;224;181;155;48;2;226;184;159m \033[38;2;223;176;149;48;2;225;182;156m \033[38;2;221;172;144;48;2;223;176;150m \033[38;2;220;172;143;48;2;222;176;147m \033[38;2;220;173;144;48;2;222;178;151m \033[38;2;216;168;137;48;2;221;176;150m \033[38;2;213;164;133;48;2;217;171;143m \033[38;2;210;163;136;48;2;214;167;138m \033[38;2;208;161;133;48;2;210;162;133m \033[38;2;205;156;129;48;2;207;156;128m \033[m");
  $display ("\033[38;2;109;84;73;48;2;104;81;64m \033[38;2;120;91;80;48;2;121;93;80m \033[38;2;121;90;78;48;2;124;90;77m \033[38;2;122;89;74;48;2;127;90;73m \033[38;2;122;88;70;48;2;128;92;73m \033[38;2;122;89;70;48;2;129;93;74m \033[38;2;122;88;72;48;2;130;94;76m \033[38;2;119;84;74;48;2;127;87;78m \033[38;2;107;74;71;48;2;119;83;81m \033[38;2;87;59;56;48;2;100;66;67m \033[38;2;75;42;44;48;2;85;49;55m \033[38;2;74;35;35;48;2;91;55;54m \033[38;2;78;39;35;48;2;111;68;62m \033[38;2;89;42;39;48;2;109;64;60m \033[38;2;100;49;49;48;2;113;65;61m \033[38;2;106;53;51;48;2;123;74;65m \033[38;2;117;65;65;48;2;141;96;91m \033[38;2;134;82;84;48;2;149;101;99m \033[38;2;143;88;89;48;2;151;99;97m \033[38;2;155;99;98;48;2;160;109;103m \033[38;2;165;113;111;48;2;176;129;125m \033[38;2;180;135;130;48;2;190;153;144m \033[38;2;191;154;148;48;2;202;174;168m \033[38;2;199;167;163;48;2;204;175;170m \033[38;2;203;169;162;48;2;212;184;172m \033[38;2;209;173;165;48;2;229;203;192m \033[38;2;223;193;185;48;2;236;207;196m \033[38;2;227;196;182;48;2;231;198;184m \033[38;2;224;183;162;48;2;225;184;162m \033[38;2;220;174;151;48;2;223;179;154m \033[38;2;220;175;151;48;2;223;178;155m \033[38;2;221;175;154;48;2;223;177;153m \033[38;2;221;174;152;48;2;221;173;144m \033[38;2;220;172;146;48;2;221;173;144m \033[38;2;218;171;143;48;2;218;171;142m \033[38;2;214;169;139;48;2;214;165;132m \033[38;2;213;165;135;48;2;211;160;129m \033[38;2;209;163;138;48;2;209;161;136m \033[38;2;206;161;134;48;2;207;161;135m \033[38;2;202;155;128;48;2;204;157;131m \033[m");
  $display ("\033[49m \033[49;38;2;117;87;79m \033[38;2;111;85;74;48;2;119;89;77m \033[38;2;113;84;73;48;2;118;87;74m \033[38;2;116;84;72;48;2;119;86;71m \033[38;2;117;83;72;48;2;120;86;71m \033[38;2;121;82;72;48;2;121;84;71m \033[38;2;120;84;76;48;2;116;81;72m \033[38;2;124;85;72;48;2;112;76;69m \033[38;2;126;85;70;48;2;108;73;64m \033[38;2;127;83;78;48;2;102;66;62m \033[38;2;124;84;76;48;2;107;70;65m \033[38;2;129;88;78;48;2;101;59;53m \033[38;2;124;78;75;48;2;85;39;37m \033[38;2;116;70;70;48;2;80;30;32m \033[38;2;100;49;53;48;2;92;38;36m \033[38;2;95;42;46;48;2;107;54;54m \033[38;2;105;50;59;48;2;121;67;70m \033[38;2;102;45;45;48;2;127;67;72m \033[38;2;97;41;37;48;2;128;62;65m \033[38;2;105;49;44;48;2;128;64;63m \033[38;2;108;53;48;48;2;140;78;73m \033[38;2;106;54;48;48;2;153;96;88m \033[38;2;110;56;52;48;2;164;114;107m \033[38;2;118;68;62;48;2;177;135;126m \033[38;2;132;86;81;48;2;180;141;128m \033[38;2;149;106;108;48;2;190;159;147m \033[38;2;176;135;133;48;2;211;177;164m \033[38;2;202;161;150;48;2;216;173;153m \033[38;2;203;160;138;48;2;214;167;143m \033[38;2;205;158;134;48;2;215;168;142m \033[38;2;208;162;141;48;2;216;168;146m \033[38;2;209;162;142;48;2;216;166;144m \033[38;2;207;160;138;48;2;214;165;141m \033[38;2;205;158;135;48;2;212;164;139m \033[38;2;202;156;130;48;2;209;162;134m \033[38;2;201;156;130;48;2;207;161;133m \033[38;2;200;155;130;48;2;206;160;134m \033[38;2;197;153;126;48;2;202;157;130m \033[38;2;196;149;124;48;2;198;151;125m \033[m");
  $display ("\033[49m  \033[49;38;2;97;73;73m \033[38;2;109;84;77;48;2;112;84;75m \033[38;2;113;86;75;48;2;114;83;73m \033[38;2;113;83;70;48;2;116;82;71m \033[38;2;115;83;69;48;2;121;86;74m \033[38;2;118;85;73;48;2;124;92;81m \033[38;2;125;90;74;48;2;131;97;80m \033[38;2;135;97;75;48;2;137;100;83m \033[38;2;150;107;93;48;2;149;105;98m \033[38;2;161;115;104;48;2;149;102;94m \033[38;2;166;124;110;48;2;146;101;89m \033[38;2;178;141;135;48;2;148;102;96m \033[38;2;168;125;123;48;2;140;92;90m \033[38;2;153;104;104;48;2;135;85;87m \033[38;2;143;90;90;48;2;131;79;82m \033[38;2;143;91;94;48;2;130;78;83m \033[38;2;147;97;97;48;2;129;79;78m \033[38;2;152;103;99;48;2;121;71;63m \033[38;2;159;107;105;48;2;120;68;65m \033[38;2;164;110;108;48;2;117;63;59m \033[38;2;169;112;112;48;2;116;57;53m \033[38;2;166;107;103;48;2;119;60;63m \033[38;2;155;100;93;48;2;115;60;67m \033[38;2;148;101;88;48;2;111;60;69m \033[38;2;142;95;76;48;2;112;64;66m \033[38;2;129;81;63;48;2;140;90;89m \033[38;2;138;90;77;48;2;169;124;116m \033[38;2;159;113;100;48;2;183;137;123m \033[38;2;173;131;114;48;2;189;143;122m \033[38;2;180;133;116;48;2;192;145;124m \033[38;2;182;134;115;48;2;194;147;125m \033[38;2;182;133;114;48;2;196;149;127m \033[38;2;183;134;114;48;2;195;149;124m \033[38;2;182;134;113;48;2;193;147;122m \033[38;2;183;136;115;48;2;193;148;123m \033[38;2;185;139;118;48;2;193;148;125m \033[38;2;186;140;122;48;2;192;147;124m \033[38;2;186;142;124;48;2;192;146;124m \033[m");
  $display ("\033[49m   \033[49;38;2;85;57;42m \033[38;2;75;60;45;48;2;104;79;65m \033[38;2;96;73;58;48;2;108;82;68m \033[38;2;103;78;66;48;2;110;80;67m \033[38;2;107;79;64;48;2;112;80;67m \033[38;2;113;80;64;48;2;116;82;64m \033[38;2;114;81;60;48;2;121;83;63m \033[38;2;116;83;60;48;2;131;88;70m \033[38;2;123;86;67;48;2;147;101;88m \033[38;2;146;97;83;48;2;163;116;106m \033[38;2;156;106;96;48;2;175;133;127m \033[38;2;166;113;107;48;2;176;132;127m \033[38;2;170;116;112;48;2;172;125;121m \033[38;2;170;115;109;48;2;168;118;117m \033[38;2;177;127;120;48;2;167;116;117m \033[38;2;194;148;144;48;2;170;122;122m \033[38;2;198;157;151;48;2;175;128;124m \033[38;2;198;157;151;48;2;180;130;126m \033[38;2;199;155;149;48;2;183;130;124m \033[38;2;199;157;146;48;2;185;133;126m \033[38;2;201;156;146;48;2;184;132;123m \033[38;2;196;152;143;48;2;178;128;117m \033[38;2;181;142;125;48;2;169;128;111m \033[38;2;176;133;117;48;2;160;116;98m \033[38;2;165;122;104;48;2;153;108;90m \033[38;2;158;115;101;48;2;143;96;82m \033[38;2;155;111;97;48;2;149;102;89m \033[38;2;158;113;101;48;2;164;118;105m \033[38;2;164;120;104;48;2;171;125;109m \033[38;2;170;125;105;48;2;175;129;109m \033[38;2;172;127;108;48;2;177;129;111m \033[38;2;173;129;110;48;2;176;130;111m \033[38;2;173;130;110;48;2;176;130;111m \033[38;2;174;130;110;48;2;177;130;113m \033[38;2;173;130;112;48;2;179;133;116m \033[38;2;172;131;113;48;2;179;136;120m \033[38;2;171;131;115;48;2;177;135;120m \033[m");
end endtask

task YOU_PASS_task; begin
    $display ("\033[38;2;15;15;16;48;2;17;15;15m \033[38;2;16;16;17;48;2;18;18;19m \033[38;2;13;13;13;48;2;15;14;15m \033[38;2;14;13;14;48;2;13;12;13m \033[38;2;14;13;14;48;2;13;13;13m \033[38;2;13;13;13;48;2;13;13;14m \033[38;2;14;14;16;48;2;14;14;15m \033[38;2;14;15;17;48;2;13;13;13m \033[38;2;16;17;18;48;2;15;15;17m \033[38;2;15;15;18;48;2;16;16;18m \033[38;2;14;15;18;48;2;14;14;16m \033[38;2;15;15;18;48;2;17;17;18m \033[38;2;17;18;21;48;2;18;18;20m \033[38;2;15;15;18;48;2;16;17;19m \033[38;2;15;15;17;48;2;17;17;19m \033[38;2;16;16;18;48;2;14;14;17m \033[38;2;12;12;17;48;2;13;12;17m \033[38;2;9;10;17;48;2;13;12;17m \033[38;2;11;11;16;48;2;13;13;17m \033[38;2;13;13;17;48;2;15;13;17m \033[38;2;15;14;18;48;2;16;14;18m \033[38;2;14;13;17;48;2;16;15;18m \033[38;2;16;14;19;48;2;18;17;20m \033[38;2;18;17;20;48;2;18;18;21m \033[38;2;18;17;20;48;2;14;14;17m \033[38;2;11;10;15;48;2;10;7;12m \033[38;2;13;11;16;48;2;15;14;18m \033[38;2;19;16;20;48;2;19;18;21m \033[38;2;16;15;19;48;2;17;15;19m \033[38;2;17;14;21;48;2;19;16;22m \033[38;2;20;19;24;48;2;24;24;26m \033[38;2;19;18;22;48;2;19;19;20m \033[38;2;17;16;21;48;2;17;15;16m \033[38;2;17;15;19;48;2;18;16;16m \033[38;2;16;15;17;48;2;16;15;15m \033[38;2;18;18;18;48;2;19;18;20m \033[38;2;20;20;21;48;2;22;22;24m \033[38;2;21;21;23;48;2;22;22;23m \033[38;2;20;20;23;48;2;19;19;23m \033[38;2;16;18;22;48;2;14;16;23m \033[m");
    $display ("\033[38;2;17;16;16;48;2;17;15;16m \033[38;2;15;16;16;48;2;16;16;17m \033[38;2;13;13;15;48;2;13;13;13m \033[38;2;13;13;16;48;2;13;13;15m \033[38;2;14;14;17;48;2;13;13;17m \033[38;2;15;16;18;48;2;13;13;15m \033[38;2;13;14;17;48;2;14;15;17m \033[38;2;13;13;16;48;2;15;15;18m \033[38;2;16;16;18;48;2;17;18;20m \033[38;2;14;14;17;48;2;13;14;16m \033[38;2;14;15;17;48;2;16;17;19m \033[38;2;13;14;16;48;2;14;14;16m \033[38;2;10;9;14;48;2;13;13;15m \033[38;2;9;9;14;48;2;14;14;17m \033[38;2;10;9;15;48;2;13;13;15m \033[38;2;7;9;16;48;2;14;15;18m \033[38;2;6;10;17;48;2;11;12;18m \033[38;2;8;12;18;48;2;8;11;18m \033[38;2;5;8;17;48;2;3;7;15m \033[38;2;5;6;14;48;2;9;8;15m \033[38;2;12;13;17;48;2;15;13;18m \033[38;2;11;11;15;48;2;14;13;18m \033[38;2;14;12;17;48;2;14;13;18m \033[38;2;20;17;23;48;2;19;15;21m \033[38;2;19;18;22;48;2;19;15;21m \033[38;2;19;18;21;48;2;17;14;19m \033[38;2;16;14;19;48;2;15;10;16m \033[38;2;14;11;17;48;2;16;13;18m \033[38;2;14;13;19;48;2;17;15;20m \033[38;2;12;12;17;48;2;16;14;20m \033[38;2;13;13;19;48;2;17;18;22m \033[38;2;14;14;18;48;2;18;18;22m \033[38;2;15;16;19;48;2;15;15;20m \033[38;2;15;14;19;48;2;14;14;19m \033[38;2;13;12;15;48;2;14;14;16m \033[38;2;14;13;16;48;2;16;14;16m \033[38;2;19;19;22;48;2;20;20;21m \033[38;2;21;20;23;48;2;21;22;23m \033[38;2;24;24;27;48;2;21;21;27m \033[38;2;21;22;27;48;2;18;20;23m \033[m");
    $display ("\033[38;2;18;18;16;48;2;17;17;16m \033[38;2;16;15;14;48;2;15;14;15m \033[38;2;13;11;14;48;2;13;13;16m \033[38;2;12;12;14;48;2;12;12;16m \033[38;2;12;11;12;48;2;13;13;16m \033[38;2;17;17;18;48;2;17;18;20m \033[38;2;15;14;17;48;2;16;17;18m \033[38;2;15;15;18;48;2;14;14;16m \033[38;2;13;12;15;48;2;14;14;17m \033[38;2;12;12;15;48;2;14;15;17m \033[38;2;12;13;16;48;2;14;14;17m \033[38;2;13;13;16;48;2;12;13;16m \033[38;2;10;10;15;48;2;12;12;15m \033[38;2;10;11;15;48;2;10;9;14m \033[38;2;8;12;16;48;2;4;6;14m \033[38;2;2;8;16;48;2;0;4;15m \033[38;2;2;7;16;48;2;5;8;16m \033[38;2;4;8;18;48;2;9;12;18m \033[38;2;3;8;19;48;2;6;10;18m \033[38;2;2;6;17;48;2;1;6;14m \033[38;2;3;10;15;48;2;6;12;15m \033[38;2;6;12;17;48;2;6;12;15m \033[38;2;3;6;13;48;2;6;8;13m \033[38;2;11;11;16;48;2;18;15;21m \033[38;2;20;18;20;48;2;21;19;24m \033[38;2;22;20;24;48;2;20;18;23m \033[38;2;17;14;20;48;2;16;14;18m \033[38;2;13;9;15;48;2;13;9;14m \033[38;2;11;8;14;48;2;12;10;15m \033[38;2;9;8;14;48;2;10;10;15m \033[38;2;8;10;18;48;2;11;11;16m \033[38;2;11;12;20;48;2;13;13;19m \033[38;2;8;11;19;48;2;13;14;21m \033[38;2;7;11;18;48;2;12;13;18m \033[38;2;8;11;17;48;2;11;11;17m \033[38;2;10;11;17;48;2;12;11;17m \033[38;2;14;13;19;48;2;17;16;21m \033[38;2;17;16;19;48;2;18;16;20m \033[38;2;24;24;29;48;2;24;22;29m \033[38;2;27;28;33;48;2;25;27;31m \033[m");
    $display ("\033[38;2;18;17;18;48;2;19;18;18m \033[38;2;16;15;17;48;2;15;15;15m \033[38;2;16;16;18;48;2;13;11;13m \033[38;2;12;13;13;48;2;12;12;11m \033[38;2;13;11;12;48;2;12;10;10m \033[38;2;13;13;14;48;2;16;15;17m \033[38;2;17;17;18;48;2;16;15;17m \033[38;2;13;13;15;48;2;14;13;15m \033[38;2;13;10;15;48;2;13;11;15m \033[38;2;13;11;16;48;2;12;11;15m \033[48;2;10;11;15m \033[38;2;11;12;16;48;2;13;14;17m \033[38;2;12;12;17;48;2;10;10;15m \033[48;2;10;10;15m \033[38;2;12;12;16;48;2;12;14;17m \033[38;2;6;10;17;48;2;4;9;16m \033[38;2;2;8;18;48;2;2;9;18m \033[48;2;3;8;18m \033[38;2;6;8;15;48;2;2;7;18m \033[38;2;8;9;14;48;2;2;6;16m \033[38;2;6;5;12;48;2;3;6;13m \033[38;2;9;7;17;48;2;9;9;17m \033[38;2;10;7;18;48;2;6;4;16m \033[38;2;8;7;17;48;2;7;8;16m \033[38;2;11;11;14;48;2;12;12;15m \033[38;2;18;16;18;48;2;21;19;23m \033[38;2;26;22;27;48;2;21;18;24m \033[38;2;13;13;23;48;2;12;9;17m \033[38;2;8;7;19;48;2;9;8;16m \033[38;2;7;6;18;48;2;6;8;16m \033[38;2;2;3;15;48;2;3;7;16m \033[38;2;1;5;14;48;2;2;6;16m \033[38;2;1;8;14;48;2;2;7;17m \033[38;2;6;11;16;48;2;5;11;18m \033[38;2;5;12;16;48;2;7;11;18m \033[38;2;6;11;15;48;2;9;11;17m \033[38;2;10;10;16;48;2;12;12;17m \033[38;2;13;12;16;48;2;15;16;18m \033[38;2;30;24;24;48;2;26;26;27m \033[38;2;36;33;33;48;2;30;32;34m \033[m");
    $display ("\033[38;2;18;17;18;48;2;18;18;18m \033[38;2;17;15;17;48;2;16;16;16m \033[38;2;17;16;18;48;2;19;19;20m \033[38;2;17;15;17;48;2;16;15;16m \033[38;2;15;14;15;48;2;14;13;12m \033[38;2;15;14;15;48;2;16;15;16m \033[38;2;13;12;12;48;2;16;15;15m \033[48;2;15;14;14m \033[38;2;13;11;15;48;2;12;9;14m \033[38;2;13;11;17;48;2;13;11;15m \033[38;2;8;9;14;48;2;7;10;14m \033[38;2;0;7;12;48;2;4;8;13m \033[38;2;1;7;12;48;2;8;10;15m \033[38;2;1;7;12;48;2;6;10;15m \033[38;2;2;4;9;48;2;9;10;15m \033[38;2;9;7;11;48;2;9;11;16m \033[38;2;9;9;13;48;2;6;9;15m \033[38;2;9;9;14;48;2;7;7;13m \033[38;2;7;7;13;48;2;5;4;11m \033[38;2;9;9;15;48;2;9;10;16m \033[38;2;16;16;21;48;2;12;13;18m \033[38;2;14;13;19;48;2;10;9;17m \033[38;2;11;9;19;48;2;10;9;19m \033[38;2;7;4;17;48;2;7;4;16m \033[38;2;10;10;19;48;2;11;11;17m \033[38;2;16;15;21;48;2;17;14;18m \033[38;2;25;22;28;48;2;28;23;27m \033[38;2;26;22;28;48;2;22;19;27m \033[38;2;8;8;18;48;2;8;7;18m \033[38;2;3;7;19;48;2;5;5;17m \033[38;2;1;7;17;48;2;1;5;15m \033[38;2;0;8;13;48;2;0;6;12m \033[48;2;0;7;12m \033[38;2;2;6;11;48;2;2;8;13m \033[38;2;5;7;13;48;2;3;9;14m \033[38;2;9;11;15;48;2;4;10;15m \033[38;2;15;13;13;48;2;11;12;13m \033[38;2;38;30;28;48;2;22;17;12m \033[38;2;52;45;41;48;2;38;29;26m \033[38;2;45;35;25;48;2;40;32;27m \033[m");
    $display ("\033[38;2;13;11;10;48;2;14;16;15m \033[38;2;17;16;18;48;2;17;15;18m \033[38;2;13;13;14;48;2;16;15;16m \033[38;2;13;13;16;48;2;15;14;16m \033[38;2;11;11;16;48;2;13;12;14m \033[38;2;12;11;14;48;2;14;13;14m \033[38;2;14;13;13;48;2;13;12;12m \033[38;2;13;12;12;48;2;13;13;12m \033[38;2;14;13;13;48;2;15;12;14m \033[38;2;17;15;18;48;2;15;13;17m \033[38;2;19;15;21;48;2;13;10;15m \033[38;2;7;5;12;48;2;2;6;11m \033[38;2;4;5;12;48;2;6;7;12m \033[38;2;9;9;14;48;2;6;9;13m \033[38;2;2;7;11;48;2;0;5;10m \033[38;2;3;7;11;48;2;6;6;10m \033[38;2;12;11;17;48;2;10;10;14m \033[38;2;19;16;22;48;2;12;11;18m \033[38;2;17;13;19;48;2;10;8;13m \033[38;2;16;13;18;48;2;12;8;15m \033[38;2;21;18;24;48;2;18;17;23m \033[38;2;31;27;38;48;2;22;20;28m \033[38;2;18;12;23;48;2;12;9;19m \033[38;2;10;9;20;48;2;8;7;19m \033[38;2;7;8;18;48;2;8;10;19m \033[38;2;10;8;18;48;2;14;11;21m \033[38;2;15;11;20;48;2;19;14;22m \033[38;2;20;18;27;48;2;23;20;25m \033[38;2;14;11;18;48;2;10;9;17m \033[38;2;10;6;15;48;2;5;8;19m \033[38;2;11;10;14;48;2;6;7;17m \033[38;2;13;12;19;48;2;7;10;16m \033[38;2;14;10;20;48;2;8;11;17m \033[38;2;32;22;29;48;2;9;8;17m \033[38;2;46;28;30;48;2;10;7;15m \033[38;2;56;35;29;48;2;15;9;15m \033[38;2;77;48;38;48;2;23;13;19m \033[38;2;129;88;66;48;2;67;48;47m \033[38;2;148;107;83;48;2;94;71;62m \033[38;2;83;57;45;48;2;56;41;33m \033[m");
    $display ("\033[38;2;15;9;3;48;2;10;5;4m \033[38;2;15;16;13;48;2;16;16;17m \033[38;2;15;16;18;48;2;12;12;18m \033[38;2;11;10;15;48;2;10;10;16m \033[38;2;11;10;14;48;2;11;11;15m \033[38;2;10;9;14;48;2;10;8;12m \033[38;2;13;12;14;48;2;15;14;15m \033[38;2;14;13;13;48;2;15;13;13m \033[38;2;16;14;15;48;2;16;13;14m \033[38;2;20;15;21;48;2;19;16;21m \033[38;2;23;19;24;48;2;22;19;25m \033[38;2;20;16;21;48;2;17;13;20m \033[38;2;17;15;20;48;2;8;10;16m \033[38;2;15;14;20;48;2;10;10;16m \033[38;2;17;14;20;48;2;10;9;14m \033[38;2;15;11;20;48;2;10;8;15m \033[38;2;15;10;18;48;2;13;11;17m \033[38;2;15;12;19;48;2;18;15;21m \033[38;2;19;16;23;48;2;21;18;22m \033[38;2;20;16;21;48;2;21;19;24m \033[38;2;27;17;23;48;2;24;14;22m \033[38;2;47;33;39;48;2;40;31;42m \033[38;2;33;22;24;48;2;24;17;25m \033[38;2;27;19;24;48;2;15;11;22m \033[38;2;30;20;26;48;2;10;9;21m \033[38;2;47;33;34;48;2;8;9;21m \033[38;2;72;52;51;48;2;18;15;24m \033[38;2;90;70;68;48;2;33;27;36m \033[38;2;79;59;57;48;2;27;18;27m \033[38;2;70;48;43;48;2;16;11;16m \033[38;2;104;73;65;48;2;27;22;27m \033[38;2;131;93;79;48;2;38;20;31m \033[38;2;149;104;83;48;2;48;20;20m \033[38;2;163;114;90;48;2;106;76;68m \033[38;2;173;120;93;48;2;123;85;70m \033[38;2;166;115;89;48;2;132;89;71m \033[38;2;173;120;95;48;2;153;99;75m \033[38;2;181;126;97;48;2;166;112;83m \033[38;2;182;130;98;48;2;167;123;87m \033[38;2;158;106;78;48;2;126;87;62m \033[m");
    $display ("\033[38;2;50;36;29;48;2;30;20;14m \033[38;2;16;12;12;48;2;13;13;10m \033[38;2;14;14;15;48;2;15;16;16m \033[38;2;17;16;16;48;2;14;14;15m \033[38;2;19;17;19;48;2;12;11;15m \033[38;2;18;16;19;48;2;10;11;15m \033[38;2;15;11;16;48;2;13;10;14m \033[38;2;15;10;15;48;2;14;11;11m \033[38;2;16;15;15;48;2;15;14;15m \033[38;2;18;14;15;48;2;16;14;16m \033[38;2;18;14;16;48;2;20;15;18m \033[38;2;15;11;15;48;2;21;16;19m \033[38;2;17;15;18;48;2;21;16;22m \033[38;2;27;19;23;48;2;17;17;21m \033[38;2;40;25;30;48;2;18;15;21m \033[38;2;68;47;49;48;2;21;13;22m \033[38;2;74;50;52;48;2;19;6;13m \033[38;2;75;47;42;48;2;13;6;6m \033[38;2;103;74;69;48;2;25;18;21m \033[38;2;98;58;50;48;2;23;12;14m \033[38;2;141;93;82;48;2;50;31;32m \033[38;2;157;110;104;48;2;83;57;56m \033[38;2;147;104;99;48;2;78;57;55m \033[38;2;153;109;96;48;2;82;58;57m \033[38;2;169;121;98;48;2;104;76;65m \033[38;2;178;126;99;48;2;136;96;78m \033[38;2;170;120;95;48;2;156;111;91m \033[38;2;146;104;81;48;2;164;118;96m \033[38;2;92;65;51;48;2;171;122;97m \033[38;2;49;34;27;48;2;168;119;94m \033[38;2;27;20;15;48;2;159;112;88m \033[38;2;17;12;9;48;2;157;111;86m \033[38;2;11;7;5;48;2;152;107;83m \033[38;2;48;35;27;48;2;164;115;89m \033[38;2;159;114;91;48;2;178;124;97m \033[38;2;195;148;116;48;2;179;126;101m \033[38;2;201;154;118;48;2;186;134;104m \033[38;2;199;151;114;48;2;190;139;106m \033[38;2;197;143;112;48;2;192;139;109m \033[38;2;186;134;105;48;2;174;124;94m \033[m");
    $display ("\033[38;2;90;55;55;48;2;73;50;48m \033[38;2;41;27;28;48;2;24;18;18m \033[38;2;48;37;35;48;2;23;20;22m \033[38;2;55;43;40;48;2;28;24;24m \033[38;2;62;48;42;48;2;34;29;26m \033[38;2;68;53;47;48;2;36;31;28m \033[38;2;66;51;48;48;2;30;22;20m \033[38;2;69;52;49;48;2;30;22;23m \033[38;2;69;51;48;48;2;37;28;28m \033[38;2;74;53;50;48;2;45;35;36m \033[38;2;77;56;56;48;2;45;37;39m \033[38;2;71;55;54;48;2;37;30;31m \033[38;2;76;58;53;48;2;43;36;35m \033[38;2;84;63;58;48;2;61;46;47m \033[38;2;95;68;63;48;2;84;60;57m \033[38;2;104;74;65;48;2;105;76;70m \033[38;2;120;84;71;48;2;125;88;85m \033[38;2;155;106;93;48;2;146;101;96m \033[38;2;181;132;125;48;2;170;123;111m \033[38;2;191;146;139;48;2;180;132;122m \033[38;2;189;146;138;48;2;187;143;133m \033[38;2;180;133;118;48;2;177;129;116m \033[38;2;179;129;106;48;2;167;119;104m \033[38;2;180;128;102;48;2;176;126;102m \033[38;2;106;75;60;48;2;178;127;101m \033[38;2;5;4;3;48;2;131;93;73m \033[38;2;0;0;0;48;2;65;46;36m \033[38;2;5;3;3;48;2;21;15;11m \033[38;2;60;43;34;48;2;3;2;1m \033[38;2;122;88;69;48;2;4;3;2m \033[38;2;156;113;92;48;2;11;8;6m \033[38;2;179;128;107;48;2;21;14;12m \033[38;2;202;153;129;48;2;32;23;19m \033[38;2;220;173;148;48;2;88;65;52m \033[38;2;227;187;156;48;2;178;137;104m \033[38;2;232;196;166;48;2;209;170;129m \033[38;2;231;198;166;48;2;214;175;136m \033[38;2;223;189;151;48;2;212;170;135m \033[38;2;205;157;122;48;2;201;149;117m \033[38;2;193;138;107;48;2;190;136;108m \033[m");
    $display ("\033[38;2;109;74;51;48;2;93;62;48m \033[38;2;79;55;44;48;2;56;40;36m \033[38;2;99;75;62;48;2;75;58;49m \033[38;2;107;78;64;48;2;87;64;54m \033[38;2;109;78;64;48;2;92;65;56m \033[38;2;102;74;60;48;2;94;67;58m \033[38;2;64;45;39;48;2;92;66;58m \033[38;2;29;20;18;48;2;91;62;55m \033[38;2;16;10;9;48;2;89;60;54m \033[38;2;12;9;8;48;2;86;59;53m \033[38;2;16;12;11;48;2;84;57;53m \033[38;2;31;21;19;48;2;91;64;58m \033[38;2;67;47;38;48;2;116;82;68m \033[38;2;106;79;66;48;2;110;82;70m \033[38;2;113;83;70;48;2;104;75;67m \033[38;2;109;74;63;48;2;107;74;63m \033[38;2;118;81;60;48;2;119;83;66m \033[38;2;148;102;79;48;2;152;102;86m \033[38;2;180;128;109;48;2;172;121;107m \033[38;2;189;139;117;48;2;185;137;124m \033[38;2;188;132;110;48;2;186;139;129m \033[38;2;185;133;121;48;2;178;131;117m \033[38;2;182;129;113;48;2;179;129;106m \033[38;2;175;126;106;48;2;165;118;96m \033[38;2;135;98;82;48;2;44;31;25m \033[38;2;134;98;78;48;2;9;7;5m \033[38;2;165;119;94;48;2;48;34;27m \033[38;2;183;130;102;48;2;126;91;70m \033[38;2;191;135;110;48;2;177;126;100m \033[38;2;207;138;119;48;2;193;138;112m \033[38;2;227;136;128;48;2;209;144;124m \033[38;2;238;113;120;48;2;223;154;138m \033[38;2;245;139;140;48;2;234;168;155m \033[38;2;244;120;129;48;2;238;161;151m \033[38;2;245;118;129;48;2;240;151;146m \033[38;2;247;147;147;48;2;243;178;164m \033[38;2;241;124;128;48;2;240;180;160m \033[38;2;234;175;148;48;2;228;190;154m \033[38;2;212;159;124;48;2;208;160;123m \033[38;2;192;139;105;48;2;192;138;106m \033[m");
    $display ("\033[38;2;140;96;68;48;2;137;94;61m \033[38;2;115;73;54;48;2;103;70;56m \033[38;2;123;88;73;48;2;115;86;70m \033[38;2;124;92;70;48;2;117;87;69m \033[38;2;100;72;55;48;2;108;77;61m \033[38;2;37;26;20;48;2;29;20;16m \033[38;2;51;36;29;48;2;2;1;1m \033[38;2;75;53;43;48;2;7;4;3m \033[38;2;89;63;53;48;2;13;9;9m \033[38;2;94;68;58;48;2;17;12;11m \033[38;2;89;64;54;48;2;14;10;9m \033[38;2;76;54;45;48;2;8;5;4m \033[38;2;56;40;32;48;2;2;1;1m \033[38;2;75;52;42;48;2;36;26;21m \033[38;2;109;77;63;48;2;104;75;62m \033[38;2;117;82;61;48;2;110;76;60m \033[38;2;155;112;81;48;2;130;91;65m \033[38;2;219;186;159;48;2;187;147;120m \033[38;2;249;243;237;48;2;236;218;209m \033[38;2;251;243;238;48;2;239;217;204m \033[38;2;246;227;215;48;2;216;165;138m \033[38;2;237;208;191;48;2;206;147;132m \033[38;2;222;175;154;48;2;199;143;124m \033[38;2;213;164;141;48;2;194;141;121m \033[38;2;205;155;136;48;2;194;141;121m \033[38;2;199;144;126;48;2;195;143;118m \033[38;2;196;141;119;48;2;188;136;110m \033[38;2;200;146;121;48;2;189;135;108m \033[38;2;213;148;130;48;2;200;135;116m \033[38;2;229;149;138;48;2;223;137;128m \033[38;2;240;99;115;48;2;239;119;126m \033[38;2;246;118;128;48;2;243;93;111m \033[38;2;247;123;131;48;2;248;126;134m \033[38;2;244;101;116;48;2;244;94;111m \033[38;2;247;133;134;48;2;247;123;131m \033[38;2;243;122;127;48;2;246;116;126m \033[38;2;239;140;133;48;2;241;115;122m \033[38;2;231;163;138;48;2;235;161;140m \033[38;2;219;165;134;48;2;216;157;127m \033[38;2;204;154;122;48;2;197;143;111m \033[m");
    $display ("\033[38;2;136;93;68;48;2;135;94;62m \033[38;2;130;86;59;48;2;124;79;56m \033[38;2;132;94;74;48;2;128;90;73m \033[38;2;139;100;77;48;2;130;96;74m \033[38;2;147;97;77;48;2;129;93;69m \033[38;2;156;94;79;48;2;125;88;70m \033[38;2;162;94;82;48;2;124;85;70m \033[38;2;169;89;84;48;2;121;82;68m \033[38;2;181;83;85;48;2;122;81;67m \033[38;2;169;92;85;48;2;124;81;67m \033[38;2;161;85;79;48;2;119;80;65m \033[38;2;140;88;73;48;2;114;79;63m \033[38;2;135;88;70;48;2;114;80;62m \033[38;2;139;93;71;48;2;122;85;67m \033[38;2;140;96;68;48;2;126;88;69m \033[38;2;161;115;79;48;2;138;97;71m \033[38;2;202;154;115;48;2;185;135;103m \033[38;2;232;197;162;48;2;225;189;152m \033[38;2;249;238;223;48;2;251;241;230m \033[38;2;253;251;249;48;2;253;249;245m \033[38;2;251;244;236;48;2;250;240;230m \033[38;2;248;234;220;48;2;248;235;224m \033[38;2;245;225;210;48;2;243;220;209m \033[38;2;237;201;179;48;2;230;188;166m \033[38;2;223;176;148;48;2;219;170;146m \033[38;2;216;164;138;48;2;208;155;132m \033[38;2;218;169;143;48;2;208;155;130m \033[38;2;226;184;162;48;2;216;169;144m \033[38;2;232;193;172;48;2;223;176;156m \033[38;2;236;199;177;48;2;231;175;157m \033[38;2;240;203;183;48;2;240;157;153m \033[38;2;240;201;182;48;2;245;168;162m \033[38;2;239;196;175;48;2;246;161;157m \033[38;2;235;186;160;48;2;243;157;148m \033[38;2;232;181;151;48;2;240;159;144m \033[38;2;230;181;150;48;2;238;164;145m \033[38;2;227;178;147;48;2;232;172;146m \033[38;2;221;170;139;48;2;225;174;142m \033[38;2;214;163;133;48;2;216;166;135m \033[38;2;207;157;126;48;2;205;152;121m \033[m");
    $display ("\033[49;38;2;128;85;71m \033[38;2;148;97;70;48;2;137;95;60m \033[38;2;157;99;70;48;2;140;97;72m \033[38;2;190;109;99;48;2;165;106;87m \033[38;2;218;94;100;48;2;186;102;95m \033[38;2;233;78;97;48;2;213;84;93m \033[38;2;228;98;108;48;2;208;97;100m \033[38;2;236;74;96;48;2;218;86;97m \033[38;2;233;105;113;48;2;223;89;101m \033[38;2;235;91;106;48;2;214;103;105m \033[38;2;231;100;107;48;2;217;83;95m \033[38;2;213;134;117;48;2;181;108;94m \033[38;2;199;139;114;48;2;162;106;84m \033[38;2;182;130;101;48;2;156;106;82m \033[38;2;162;109;77;48;2;153;105;77m \033[38;2;164;115;78;48;2;165;118;80m \033[38;2;216;184;146;48;2;203;158;116m \033[38;2;245;224;205;48;2;243;214;189m \033[38;2;249;237;224;48;2;250;240;227m \033[38;2;252;246;238;48;2;254;253;251m \033[38;2;253;247;244;48;2;254;249;244m \033[38;2;251;240;234;48;2;251;240;232m \033[38;2;249;232;221;48;2;247;230;215m \033[38;2;246;226;214;48;2;241;213;195m \033[38;2;236;198;179;48;2;226;174;144m \033[38;2;216;160;133;48;2;217;165;138m \033[38;2;226;180;154;48;2;224;177;150m \033[38;2;234;195;174;48;2;233;192;169m \033[38;2;239;204;182;48;2;237;201;179m \033[38;2;239;207;186;48;2;240;207;185m \033[38;2;239;203;180;48;2;240;206;184m \033[38;2;236;198;170;48;2;239;203;177m \033[38;2;235;197;168;48;2;237;201;173m \033[38;2;234;195;167;48;2;233;194;165m \033[38;2;230;188;156;48;2;231;186;156m \033[38;2;227;181;149;48;2;228;182;150m \033[38;2;223;175;144;48;2;224;175;145m \033[38;2;218;169;139;48;2;219;166;137m \033[38;2;213;164;138;48;2;214;163;135m \033[38;2;209;163;137;48;2;210;163;136m \033[m");
    $display ("\033[49m \033[38;2;143;92;71;48;2;150;98;82m \033[38;2;158;107;81;48;2;171;108;87m \033[38;2;168;111;89;48;2;190;107;97m \033[38;2;185;101;91;48;2;224;80;94m \033[38;2;190;108;98;48;2;222;97;104m \033[38;2;202;111;104;48;2;229;93;105m \033[38;2;211;115;107;48;2;232;89;104m \033[38;2;217;125;115;48;2;232;112;117m \033[38;2;220;137;121;48;2;234;102;110m \033[38;2;218;153;126;48;2;228;130;120m \033[38;2;217;164;130;48;2;220;150;126m \033[38;2;217;170;132;48;2;214;159;129m \033[38;2;206;158;124;48;2;198;146;115m \033[38;2;172;114;80;48;2;159;98;64m \033[38;2;199;158;128;48;2;177;130;97m \033[38;2;207;171;134;48;2;224;201;172m \033[38;2;229;191;158;48;2;241;218;194m \033[38;2;237;202;176;48;2;245;225;207m \033[38;2;239;210;191;48;2;246;228;211m \033[38;2;233;201;179;48;2;248;233;219m \033[38;2;212;160;139;48;2;246;226;210m \033[38;2;144;99;85;48;2;242;207;191m \033[38;2;136;99;89;48;2;241;210;192m \033[38;2;218;173;144;48;2;245;221;201m \033[38;2;232;188;150;48;2;227;181;153m \033[38;2;231;189;161;48;2;227;182;158m \033[38;2;235;197;172;48;2;234;197;173m \033[38;2;236;201;174;48;2;237;202;177m \033[38;2;236;198;172;48;2;238;204;179m \033[38;2;235;192;166;48;2;237;198;173m \033[38;2;233;188;161;48;2;234;192;161m \033[38;2;232;189;159;48;2;233;191;160m \033[38;2;229;186;154;48;2;231;186;155m \033[38;2;227;183;148;48;2;227;180;145m \033[38;2;224;178;148;48;2;225;177;146m \033[38;2;222;177;149;48;2;222;177;148m \033[38;2;219;174;143;48;2;220;173;143m \033[38;2;213;164;135;48;2;214;164;137m \033[38;2;208;159;133;48;2;209;160;133m \033[m");
    $display ("\033[49m \033[38;2;128;91;55;48;2;128;89;64m \033[38;2;138;95;73;48;2;146;104;76m \033[38;2;148;111;85;48;2;152;113;82m \033[38;2;147;108;84;48;2;154;109;83m \033[38;2;155;115;86;48;2;162;113;88m \033[38;2;167;123;97;48;2;174;120;98m \033[38;2;181;132;107;48;2;186;127;104m \033[38;2;194;145;119;48;2;199;140;115m \033[38;2;204;151;123;48;2;209;150;122m \033[38;2;211;157;123;48;2;214;159;125m \033[38;2;217;166;129;48;2;218;168;130m \033[38;2;220;173;138;48;2;220;172;135m \033[38;2;217;172;139;48;2;212;165;130m \033[38;2;200;145;114;48;2;202;151;121m \033[38;2;152;99;74;48;2;191;142;116m \033[38;2;81;38;26;48;2;151;104;79m \033[38;2;80;40;30;48;2;156;116;96m \033[38;2;127;80;59;48;2;184;131;112m \033[38;2;154;104;83;48;2;195;137;113m \033[38;2;160;108;91;48;2;184;123;102m \033[38;2;159;108;91;48;2;149;96;82m \033[38;2;160;110;94;48;2;79;46;42m \033[38;2;169;114;103;48;2;65;38;34m \033[38;2;181;122;112;48;2;149;92;74m \033[38;2;190;123;108;48;2;210;149;122m \033[38;2;228;188;169;48;2;232;195;171m \033[38;2;243;220;208;48;2;237;209;185m \033[38;2;238;205;188;48;2;235;199;174m \033[38;2;221;178;156;48;2;230;190;164m \033[38;2;203;155;134;48;2;226;181;157m \033[38;2;202;152;132;48;2;223;177;153m \033[38;2;206;155;133;48;2;222;175;151m \033[38;2;208;159;134;48;2;222;175;149m \033[38;2;210;160;135;48;2;221;175;145m \033[38;2;211;163;136;48;2;220;174;145m \033[38;2;211;164;136;48;2;219;173;144m \033[38;2;211;163;137;48;2;216;170;140m \033[38;2;208;160;135;48;2;212;164;135m \033[38;2;206;159;136;48;2;207;160;135m \033[m");
    $display ("\033[49m  \033[49;38;2;134;85;73m \033[38;2;146;119;89;48;2;149;115;90m \033[38;2;146;116;92;48;2;144;108;86m \033[38;2;152;119;94;48;2;152;114;87m \033[38;2;163;124;97;48;2;164;123;95m \033[38;2;173;128;104;48;2;175;130;105m \033[38;2;180;132;108;48;2;186;138;115m \033[38;2;186;135;109;48;2;196;144;119m \033[38;2;195;139;112;48;2;204;149;119m \033[38;2;205;148;116;48;2;212;158;126m \033[38;2;212;158;123;48;2;218;169;135m \033[38;2;216;167;139;48;2;220;172;145m \033[38;2;191;137;120;48;2;181;126;102m \033[38;2;127;73;58;48;2;123;72;52m \033[38;2;121;79;67;48;2;110;72;60m \033[38;2;130;90;84;48;2;115;80;74m \033[38;2;148;107;94;48;2;134;94;75m \033[38;2;157;114;105;48;2;150;107;95m \033[38;2;154;109;99;48;2;152;109;95m \033[38;2;152;103;92;48;2;157;110;93m \033[38;2;170;121;113;48;2;170;122;104m \033[38;2;191;147;136;48;2;177;131;114m \033[38;2;205;169;159;48;2;185;141;127m \033[38;2;212;180;175;48;2;194;145;131m \033[38;2;218;189;181;48;2;224;190;174m \033[38;2;213;177;168;48;2;238;213;204m \033[38;2;182;140;134;48;2;224;193;183m \033[38;2;151;100;94;48;2;192;145;135m \033[38;2;154;102;88;48;2;168;118;104m \033[38;2;168;118;104;48;2;180;129;114m \033[38;2;179;129;113;48;2;190;139;120m \033[38;2;188;138;117;48;2;195;144;122m \033[38;2;191;141;120;48;2;197;146;124m \033[38;2;193;142;121;48;2;199;148;125m \033[38;2;193;143;121;48;2;200;150;126m \033[38;2;194;144;122;48;2;202;152;129m \033[38;2;194;146;127;48;2;201;153;132m \033[38;2;192;147;130;48;2;199;153;134m \033[m");
    $display ("\033[49m   \033[38;2;148;121;94;48;2;149;123;98m \033[38;2;144;119;93;48;2;148;121;96m \033[38;2;144;116;91;48;2;149;121;96m \033[38;2;148;114;89;48;2;158;125;97m \033[38;2;155;114;86;48;2;166;126;99m \033[38;2;161;114;87;48;2;171;124;99m \033[38;2;164;113;87;48;2;177;123;98m \033[38;2;170;116;90;48;2;183;127;100m \033[38;2;173;121;93;48;2;195;135;105m \033[38;2;170;121;94;48;2;200;141;107m \033[38;2;165;122;96;48;2;200;151;121m \033[38;2;143;103;82;48;2;192;149;128m \033[38;2;131;92;81;48;2;169;122;105m \033[38;2;133;93;87;48;2;154;113;98m \033[38;2;124;85;77;48;2;145;104;95m \033[38;2;117;71;65;48;2;147;105;94m \033[38;2;128;81;77;48;2;157;110;103m \033[38;2;135;85;85;48;2;158;105;103m \033[38;2;139;84;85;48;2;153;97;93m \033[38;2;150;88;89;48;2;170;113;109m \033[38;2;144;84;82;48;2;195;147;142m \033[38;2;142;85;79;48;2;206;165;157m \033[38;2;130;76;67;48;2;206;166;162m \033[38;2;116;63;57;48;2;192;148;141m \033[38;2;111;57;57;48;2;168;120;110m \033[38;2;120;66;70;48;2;124;72;73m \033[38;2;152;102;89;48;2;130;79;69m \033[38;2;176;129;107;48;2;166;116;97m \033[38;2;182;137;118;48;2;173;127;110m \033[38;2;177;130;114;48;2;173;125;111m \033[38;2;177;128;111;48;2;180;132;113m \033[38;2;181;133;112;48;2;187;137;118m \033[38;2;185;137;116;48;2;189;140;120m \033[38;2;186;139;117;48;2;189;140;120m \033[38;2;186;140;117;48;2;189;142;120m \033[38;2;184;139;117;48;2;189;142;121m \033[38;2;180;139;119;48;2;186;142;123m \033[m");
    $display ("\033[49m    \033[38;2;130;103;81;48;2;136;117;89m \033[38;2;130;107;85;48;2;137;111;87m \033[38;2;136;105;85;48;2;142;109;85m \033[38;2;136;104;80;48;2;148;107;82m \033[38;2;141;103;77;48;2;153;109;83m \033[38;2;143;102;76;48;2;156;109;83m \033[38;2;140;99;76;48;2;155;109;83m \033[38;2;131;94;75;48;2;148;107;81m \033[38;2;115;81;74;48;2;143;106;83m \033[38;2;91;64;65;48;2;116;85;76m \033[38;2;70;48;47;48;2;85;56;58m \033[38;2;67;40;40;48;2;72;41;43m \033[38;2;70;39;35;48;2;83;50;47m \033[38;2;71;34;28;48;2;90;52;49m \033[38;2;75;37;34;48;2;94;52;50m \033[38;2;80;40;37;48;2;97;52;50m \033[38;2;86;44;40;48;2;102;57;56m \033[38;2;95;54;54;48;2;111;62;65m \033[38;2;99;57;50;48;2;107;53;54m \033[38;2;104;63;52;48;2;95;46;41m \033[38;2;122;78;69;48;2;94;48;42m \033[38;2;144;93;84;48;2;96;49;42m \033[38;2;161;106;97;48;2;117;61;58m \033[38;2;173;117;104;48;2;140;81;81m \033[38;2;181;130;113;48;2;160;105;96m \033[38;2;187;142;124;48;2;174;129;110m \033[38;2;194;154;137;48;2;187;142;124m \033[38;2;192;152;137;48;2;191;147;130m \033[38;2;180;137;121;48;2;180;134;117m \033[38;2;174;128;109;48;2;175;127;110m \033[38;2;172;125;106;48;2;175;128;108m \033[38;2;171;125;104;48;2;177;131;109m \033[38;2;170;125;103;48;2;180;133;110m \033[38;2;172;126;104;48;2;182;135;114m \033[38;2;172;127;107;48;2;179;134;112m \033[38;2;161;121;100;48;2;176;138;115m \033[m");
    $display ("\033[49m     \033[49;38;2;121;98;80m \033[38;2;108;86;68;48;2;126;102;84m \033[38;2;129;100;86;48;2;131;98;80m \033[38;2;123;92;78;48;2;131;95;74m \033[38;2;120;87;72;48;2;130;94;72m \033[38;2;116;84;67;48;2;126;90;71m \033[38;2;112;81;66;48;2;116;85;69m \033[38;2;110;76;67;48;2;108;78;67m \033[38;2;106;73;65;48;2;96;69;63m \033[38;2;110;78;62;48;2;93;63;57m \033[38;2;114;78;65;48;2;95;64;59m \033[38;2;117;79;68;48;2;101;70;61m \033[38;2;115;80;64;48;2;102;71;59m \033[38;2;119;84;68;48;2;102;67;59m \033[38;2;122;86;71;48;2;106;68;61m \033[38;2;121;83;69;48;2;110;70;63m \033[38;2;123;84;70;48;2;115;74;66m \033[38;2;124;87;73;48;2;122;82;72m \033[38;2;133;95;78;48;2;127;87;72m \033[38;2;141;102;84;48;2;138;95;82m \033[38;2;146;106;88;48;2;149;103;87m \033[38;2;152;112;94;48;2;157;112;95m \033[38;2;160;118;101;48;2;169;124;107m \033[38;2;169;124;106;48;2;180;136;119m \033[38;2;170;128;112;48;2;188;145;127m \033[38;2;171;127;113;48;2;190;149;134m \033[38;2;169;126;112;48;2;184;143;130m \033[38;2;169;126;108;48;2;176;135;116m \033[38;2;169;123;105;48;2;173;127;108m \033[38;2;168;120;102;48;2;170;123;105m \033[38;2;163;118;99;48;2;166;120;100m \033[38;2;159;115;96;48;2;164;118;98m \033[38;2;157;114;96;48;2;163;118;96m \033[38;2;150;111;92;48;2;161;119;100m \033[38;2;131;100;77;48;2;146;109;91m \033[m");
    $display ("\033[49m      \033[49;38;2;73;55;36m \033[49;38;2;108;84;70m \033[38;2;109;84;73;48;2;125;94;85m \033[38;2;114;90;76;48;2;116;87;74m \033[38;2;112;84;72;48;2;114;83;70m \033[38;2;110;80;69;48;2;112;81;69m \033[38;2;113;81;70;48;2;111;77;68m \033[38;2;116;86;72;48;2;114;82;71m \033[38;2;118;86;69;48;2;118;85;70m \033[38;2;119;86;66;48;2;120;87;70m \033[38;2;122;86;67;48;2;125;88;72m \033[38;2;124;87;68;48;2;124;87;70m \033[38;2;127;89;72;48;2;126;91;73m \033[38;2;129;90;73;48;2;129;94;77m \033[38;2;130;91;73;48;2;126;91;74m \033[38;2;132;91;73;48;2;128;90;73m \033[38;2;135;95;74;48;2;129;91;73m \033[38;2;139;97;79;48;2;137;98;80m \033[38;2;143;98;80;48;2;141;101;83m \033[38;2;143;101;82;48;2;143;103;84m \033[38;2;145;100;83;48;2;146;105;87m \033[38;2;146;103;83;48;2;148;105;87m \033[38;2;150;106;88;48;2;151;107;89m \033[38;2;154;110;94;48;2;154;111;94m \033[38;2;157;115;98;48;2;158;113;97m \033[38;2;158;115;100;48;2;159;115;98m \033[38;2;156;112;98;48;2;162;117;100m \033[38;2;154;112;97;48;2;161;117;101m \033[38;2;153;113;95;48;2;161;115;99m \033[38;2;150;113;94;48;2;158;114;98m \033[38;2;143;109;93;48;2;153;113;95m \033[38;2;139;107;90;48;2;148;110;94m \033[49;38;2;145;106;89m \033[49m \033[m");

    $display ("--------------------------------------------------------------------");
    $display ("                  You have passed all patterns!                     ");
    $display ("                  Total latency : %d cycles                     ", total_latency);
    $display ("--------------------------------------------------------------------");
end endtask


endprogram